magic
tech sky130A
magscale 1 2
timestamp 1731032193
<< locali >>
rect 2884 5173 4988 5188
rect 2884 5126 3030 5173
rect 4872 5126 4988 5173
rect 2884 5112 4988 5126
rect 2884 5095 2960 5112
rect 1160 4840 2668 4850
rect 1160 4780 1186 4840
rect 1148 4770 1186 4780
rect 2646 4780 2668 4840
rect 2646 4770 2682 4780
rect 1148 4713 2682 4770
rect 1148 4704 2621 4713
rect 548 3690 624 3694
rect 1148 3690 1224 4704
rect 1887 4644 1949 4704
rect 548 3650 1224 3690
rect 548 930 560 3650
rect 615 3614 1224 3650
rect 615 930 624 3614
rect 548 378 624 930
rect 1149 3469 1224 3614
rect 1149 378 1162 3469
rect 548 334 1162 378
rect 1205 378 1224 3469
rect 1888 4630 1949 4644
rect 1888 378 1897 4630
rect 1205 351 1897 378
rect 1943 378 1949 4630
rect 2606 751 2621 4704
rect 2669 751 2682 4713
rect 2606 378 2682 751
rect 1943 351 2682 378
rect 1205 334 2682 351
rect 548 302 2682 334
rect 2884 700 2901 5095
rect 2941 700 2960 5095
rect 1149 301 1224 302
rect 514 74 2794 142
rect 514 -1226 582 74
rect 1252 -1226 1323 74
rect 1994 -1226 2060 74
rect 2726 -1226 2794 74
rect 514 -1242 2794 -1226
rect 514 -1302 576 -1242
rect 2750 -1302 2794 -1242
rect 514 -1308 2794 -1302
rect 530 -1310 2794 -1308
rect 2884 -1226 2960 700
rect 4912 5091 4988 5112
rect 4912 -1197 4927 5091
rect 4978 -1197 4988 5091
rect 4912 -1226 4988 -1197
rect 2884 -1242 4988 -1226
rect 2884 -1294 2946 -1242
rect 4950 -1258 4988 -1242
rect 4950 -1294 4990 -1258
rect 530 -1316 2774 -1310
rect 2884 -1334 4990 -1294
<< viali >>
rect 3030 5126 4872 5173
rect 1186 4770 2646 4840
rect 560 930 615 3650
rect 1162 334 1205 3469
rect 1897 351 1943 4630
rect 2621 751 2669 4713
rect 2901 700 2941 5095
rect 576 -1302 2750 -1242
rect 4927 -1197 4978 5091
rect 2946 -1294 4950 -1242
<< metal1 >>
rect 2886 5189 4987 5191
rect 1632 5150 2004 5178
rect 1632 4850 1664 5150
rect 1160 4840 1664 4850
rect 1972 4850 2004 5150
rect 2885 5173 4987 5189
rect 2885 5126 3030 5173
rect 4872 5126 4987 5173
rect 2885 5112 4987 5126
rect 2885 5095 2960 5112
rect 2610 4850 2683 4851
rect 1972 4842 2683 4850
rect 1972 4840 2052 4842
rect 1160 4770 1186 4840
rect 2648 4772 2683 4842
rect 2646 4770 2683 4772
rect 1160 4713 2683 4770
rect 1160 4710 2621 4713
rect 1145 4582 1746 4636
rect 1145 4576 1384 4582
rect 549 3650 626 3695
rect 549 930 560 3650
rect 615 930 626 3650
rect 1145 3587 1199 4576
rect 785 3533 1199 3587
rect 1256 4122 1310 4534
rect 1149 3469 1224 3492
rect 724 1698 1040 2090
rect 549 902 626 930
rect 701 486 747 502
rect 1029 486 1075 502
rect 701 444 1075 486
rect 482 52 682 178
rect 858 52 954 444
rect 1149 334 1162 3469
rect 1205 334 1224 3469
rect 1149 301 1224 334
rect 1256 477 1320 4122
rect 1502 330 1598 4582
rect 1780 534 1850 4710
rect 1888 4630 1949 4658
rect 1256 240 1320 326
rect 1158 176 1320 240
rect 1496 310 1598 330
rect 1888 351 1897 4630
rect 1943 351 1949 4630
rect 1496 298 1806 310
rect 1888 302 1949 351
rect 1990 312 2038 4522
rect 2228 494 2324 4632
rect 2501 621 2547 4525
rect 2610 751 2621 4710
rect 2669 751 2683 4713
rect 2610 733 2683 751
rect 2885 700 2901 5095
rect 2941 700 2960 5095
rect 4912 5091 4987 5112
rect 3048 4616 3708 5050
rect 3804 4616 4464 5050
rect 2885 677 2960 700
rect 2495 592 2874 621
rect 2495 575 2784 592
rect 2184 430 2377 494
rect 2184 366 2190 430
rect 2371 366 2377 430
rect 1496 240 1518 298
rect 1790 240 1806 298
rect 1990 264 2680 312
rect 1496 234 1806 240
rect 1500 228 1806 234
rect 2118 188 2448 198
rect 482 -22 1112 52
rect 550 -660 678 -88
rect 550 -1226 558 -660
rect 530 -1278 558 -1226
rect 858 -1122 954 -22
rect 1158 -94 1222 176
rect 2118 134 2126 188
rect 2438 134 2448 188
rect 2118 124 2448 134
rect 1110 -572 1222 -94
rect 1292 -666 1420 -88
rect 1292 -1064 1298 -666
rect 1292 -1080 1420 -1064
rect 1608 -1122 1704 -58
rect 1878 -476 1924 -102
rect 2126 -476 2174 -88
rect 1878 -674 2174 -476
rect 1878 -1086 1924 -674
rect 1864 -1122 1924 -1086
rect 2126 -1096 2174 -674
rect 720 -1178 1924 -1122
rect 2352 -1158 2448 124
rect 2632 -1078 2680 264
rect 2772 242 2784 575
rect 2856 242 2874 592
rect 2772 228 2874 242
rect 2828 -750 2874 228
rect 722 -1192 1924 -1178
rect 2828 -1182 3330 -750
rect 3426 -1184 4086 -750
rect 4180 -1184 4840 -750
rect 4912 -1197 4927 5091
rect 4978 -1197 4987 5091
rect 4912 -1226 4987 -1197
rect 680 -1242 2774 -1226
rect 530 -1302 576 -1278
rect 2750 -1302 2774 -1242
rect 530 -1316 2774 -1302
rect 2916 -1242 4987 -1226
rect 2916 -1294 2946 -1242
rect 4950 -1294 4987 -1242
rect 2916 -1312 4987 -1294
rect 4912 -1316 4987 -1312
<< via1 >>
rect 1664 4840 1972 5150
rect 2052 4840 2648 4842
rect 1186 4770 1606 4840
rect 1664 4832 1972 4840
rect 2052 4772 2646 4840
rect 2646 4772 2648 4840
rect 1256 326 1320 477
rect 4577 4634 4827 5031
rect 2190 366 2371 430
rect 1518 240 1790 298
rect 558 -1242 680 -660
rect 2126 134 2438 188
rect 1298 -1064 1420 -666
rect 2784 242 2856 592
rect 558 -1278 576 -1242
rect 576 -1278 680 -1242
rect 762 -1296 2736 -1244
rect 2946 -1294 4950 -1242
<< metal2 >>
rect 1069 5150 5039 5225
rect 1069 4840 1664 5150
rect 1069 4770 1186 4840
rect 1606 4832 1664 4840
rect 1972 5031 5039 5150
rect 1972 4842 4577 5031
rect 1972 4832 2052 4842
rect 1606 4772 2052 4832
rect 2648 4772 4577 4842
rect 1606 4770 4577 4772
rect 1069 4634 4577 4770
rect 4827 4634 5039 5031
rect 1069 4517 5039 4634
rect 2772 592 2870 608
rect 1256 477 1320 484
rect 511 190 679 327
rect 1320 366 2190 430
rect 2371 366 2377 430
rect 1256 319 1320 326
rect 2772 310 2784 592
rect 1500 298 2784 310
rect 1500 240 1518 298
rect 1790 242 2784 298
rect 2856 242 2870 592
rect 1790 240 2870 242
rect 1500 228 2870 240
rect 2118 190 2448 198
rect 511 188 2459 190
rect 511 134 2126 188
rect 2438 134 2459 188
rect 511 128 2459 134
rect 511 127 679 128
rect 2118 124 2448 128
rect 323 -660 5033 -639
rect 323 -1278 558 -660
rect 680 -666 5033 -660
rect 680 -1064 1298 -666
rect 1420 -1064 5033 -666
rect 680 -1242 5033 -1064
rect 680 -1244 2946 -1242
rect 680 -1278 762 -1244
rect 323 -1296 762 -1278
rect 2736 -1294 2946 -1244
rect 4950 -1294 5033 -1242
rect 2736 -1296 5033 -1294
rect 323 -1347 5033 -1296
use sky130_fd_pr__nfet_g5v0d10v5_35MXHD  XM1 paramcells
timestamp 1731019923
transform 1 0 913 0 1 -591
box -436 -758 436 758
use sky130_fd_pr__nfet_g5v0d10v5_35MXHD  XM2
timestamp 1731019923
transform 1 0 1655 0 1 -591
box -436 -758 436 758
use sky130_fd_pr__pfet_g5v0d10v5_VXYCT5  XM3 paramcells
timestamp 1731019923
transform 1 0 1553 0 1 2535
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_VXYCT5  XM4
timestamp 1731019923
transform 1 0 2279 0 1 2535
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_G59KN9  XM5 paramcells
timestamp 1731019923
transform 0 1 888 -1 0 1996
box -1758 -397 1758 397
use sky130_fd_pr__nfet_g5v0d10v5_35MXHD  XM8
timestamp 1731019923
transform 1 0 2397 0 1 -591
box -436 -758 436 758
use sky130_fd_pr__res_high_po_1p41_3L9D94  XR2 paramcells
timestamp 1731019923
transform -1 0 3946 0 -1 1933
box -1063 -3282 1063 3282
<< labels >>
flabel metal2 2529 4975 2729 5175 0 FreeSans 256 90 0 0 VDD
port 0 nsew
flabel metal2 4794 -1104 4994 -904 0 FreeSans 256 90 0 0 VSS
port 1 nsew
flabel metal1 482 -22 682 178 0 FreeSans 256 90 0 0 VBN
port 2 nsew
flabel metal2 511 127 679 327 0 FreeSans 256 90 0 0 ena3v3
port 3 nsew
<< end >>
