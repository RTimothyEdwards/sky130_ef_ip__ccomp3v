magic
tech sky130A
magscale 1 2
timestamp 1717782065
<< error_s >>
rect 10123 2291 10124 4242
rect 1475 -2520 3259 -2516
rect 3257 -2566 3259 -2520
rect 1497 -2601 3237 -2595
rect 1497 -2635 3237 -2629
rect 3229 -2690 3231 -2662
rect 1503 -2716 3231 -2715
rect 3257 -2716 3259 -2690
<< dnwell >>
rect -91 -2456 11101 10125
<< nwell >>
rect -200 10017 11210 10234
rect -200 -2250 115 10017
rect 10377 6187 11210 10017
rect 5141 5929 11210 6187
rect 9361 5860 11210 5929
rect 10895 -2250 11210 5860
rect -200 -2565 11210 -2250
<< mvpsubdiff >>
rect -322 10323 -262 10357
rect 11277 10323 11337 10357
rect -322 10297 -288 10323
rect 11303 10297 11337 10323
rect -322 -2656 -288 -2630
rect 11303 -2656 11337 -2630
rect -322 -2690 -262 -2656
rect 11277 -2690 11337 -2656
<< mvnsubdiff >>
rect -134 10148 11144 10168
rect -134 10114 -54 10148
rect 11064 10114 11144 10148
rect -134 10094 11144 10114
rect -134 10088 -60 10094
rect -134 -2419 -114 10088
rect -80 -2419 -60 10088
rect -134 -2425 -60 -2419
rect 11070 10088 11144 10094
rect 11070 5833 11090 10088
rect 11124 5833 11144 10088
rect 11070 5785 11144 5833
rect 11070 5730 11090 5785
rect 11124 5730 11144 5785
rect 11070 5575 11144 5730
rect 11070 -2410 11090 5575
rect 11124 -2410 11144 5575
rect 11070 -2425 11144 -2410
rect -134 -2445 11144 -2425
rect -134 -2479 -54 -2445
rect 11054 -2479 11144 -2445
rect -134 -2499 11144 -2479
<< mvpsubdiffcont >>
rect -262 10323 11277 10357
rect -322 -2630 -288 10297
rect 11303 -2630 11337 10297
rect -262 -2690 11277 -2656
<< mvnsubdiffcont >>
rect -54 10114 11064 10148
rect -114 -2419 -80 10088
rect 11090 5833 11124 10088
rect 11090 5730 11124 5785
rect 11090 -2410 11124 5575
rect -54 -2479 11054 -2445
<< locali >>
rect -322 10323 -262 10357
rect 11277 10323 11337 10357
rect -322 10317 11337 10323
rect -322 10297 -180 10317
rect -288 10268 -180 10297
rect 11175 10297 11337 10317
rect 11175 10268 11303 10297
rect -288 10235 11303 10268
rect -288 10154 -201 10235
rect -288 -2490 -276 10154
rect -224 -2490 -201 10154
rect 11209 10193 11303 10235
rect -114 10114 -54 10148
rect 11064 10114 11124 10148
rect -114 10088 11124 10114
rect -80 10065 11090 10088
rect -80 10015 84 10065
rect 10905 10015 11090 10065
rect -80 9970 11090 10015
rect -80 9936 63 9970
rect -80 -2285 -59 9936
rect -5 -2285 63 9936
rect 10935 9915 11090 9970
rect 10935 5851 10980 9915
rect 11032 5851 11090 9915
rect 10935 5833 11090 5851
rect -80 -2290 63 -2285
rect 10934 5785 11124 5833
rect 10934 5730 11090 5785
rect 10934 5713 11124 5730
rect 10934 -2290 10980 5713
rect -80 -2297 10980 -2290
rect 11036 5575 11124 5713
rect 11036 -2297 11090 5575
rect -80 -2352 11090 -2297
rect -80 -2405 32 -2352
rect 10929 -2405 11090 -2352
rect -80 -2410 11090 -2405
rect -80 -2419 11124 -2410
rect -114 -2445 11124 -2419
rect -114 -2479 -54 -2445
rect 11054 -2479 11124 -2445
rect -288 -2566 -201 -2490
rect 11209 -2538 11237 10193
rect 11294 -2538 11303 10193
rect 11209 -2566 11303 -2538
rect -288 -2595 11303 -2566
rect -288 -2630 -153 -2595
rect -322 -2635 -153 -2630
rect 11184 -2630 11303 -2595
rect 11184 -2635 11337 -2630
rect -322 -2656 11337 -2635
rect -322 -2690 -262 -2656
rect 11277 -2690 11337 -2656
<< viali >>
rect -180 10268 11175 10317
rect -276 -2490 -224 10154
rect 84 10015 10905 10065
rect -59 -2285 -5 9936
rect 10980 5851 11032 9915
rect 10980 -2297 11036 5713
rect 32 -2405 10929 -2352
rect 11237 -2538 11294 10193
rect -153 -2635 11184 -2595
<< metal1 >>
rect -322 10317 11337 10357
rect -322 10268 -180 10317
rect 11175 10268 11337 10317
rect -322 10235 11337 10268
rect -322 10154 -201 10235
rect -322 -2490 -276 10154
rect -224 -2490 -201 10154
rect 11209 10193 11337 10235
rect -72 10065 11050 10085
rect -72 10015 84 10065
rect 10905 10015 11050 10065
rect -72 10002 11050 10015
rect -72 9936 11 10002
rect 5161 9987 5347 10002
rect -72 -2285 -59 9936
rect -5 -2285 11 9936
rect 10967 9915 11050 10002
rect 10967 6175 10980 9915
rect 10866 6164 10980 6175
rect 11032 6175 11050 9915
rect 11209 7635 11237 10193
rect 11137 7627 11237 7635
rect 11294 7627 11337 10193
rect 11032 6164 11072 6175
rect 10866 5944 10875 6164
rect 11061 5944 11072 6164
rect 10866 5935 10980 5944
rect -72 -2334 11 -2285
rect 10967 5851 10980 5935
rect 11032 5936 11072 5944
rect 11032 5935 11063 5936
rect 11032 5851 11050 5935
rect 11309 5899 11337 7627
rect 11137 5891 11237 5899
rect 10967 5713 11050 5851
rect 10967 -2297 10980 5713
rect 11036 -2297 11050 5713
rect 10967 -2334 11050 -2297
rect -72 -2352 11050 -2334
rect -72 -2405 32 -2352
rect 10929 -2405 11050 -2352
rect -72 -2417 11050 -2405
rect -322 -2520 -201 -2490
rect -322 -2544 3257 -2520
rect -322 -2595 1503 -2544
rect 3231 -2566 3257 -2544
rect 11209 -2538 11237 5891
rect 11294 -2538 11337 5899
rect 11209 -2566 11337 -2538
rect 3231 -2595 11337 -2566
rect -322 -2635 -153 -2595
rect 11184 -2635 11337 -2595
rect -322 -2690 1503 -2635
rect -319 -2716 1503 -2690
rect 3231 -2690 11337 -2635
rect 3231 -2716 3257 -2690
rect -319 -2743 3257 -2716
<< via1 >>
rect 10875 5944 10980 6164
rect 10980 5944 11032 6164
rect 11032 5944 11061 6164
rect 11137 5899 11237 7627
rect 11237 5899 11294 7627
rect 11294 5899 11309 7627
<< metal2 >>
rect 5161 9987 5347 10085
rect 11113 7627 11336 7653
rect 4961 6175 5147 6257
rect 9712 6164 11072 6175
rect 9712 6163 10875 6164
rect 9712 5949 9725 6163
rect 10824 5949 10875 6163
rect 9712 5944 10875 5949
rect 11061 5944 11072 6164
rect 9712 5936 11072 5944
rect 9712 5935 11063 5936
rect 4961 5914 5147 5935
rect 11113 5899 11137 7627
rect 11309 5899 11336 7627
rect 11113 4077 11336 5899
rect 10640 3417 11337 3922
rect -140 1871 198 1971
rect 10897 1738 11337 1838
rect -140 1636 198 1736
<< via2 >>
rect 4961 5935 5147 6175
rect 9725 5949 10824 6163
<< metal3 >>
rect 623 2142 723 7084
rect 1659 6114 1759 7545
rect 4954 6175 5158 6184
rect 835 6014 1759 6114
rect 2077 6160 4961 6175
rect 835 1343 935 6014
rect 2077 5948 2090 6160
rect 2488 5948 4961 6160
rect 2077 5935 4961 5948
rect 5147 6163 11014 6175
rect 5147 5949 9725 6163
rect 10824 5949 11014 6163
rect 5147 5935 11014 5949
rect 4954 5927 5158 5935
<< via3 >>
rect 2090 5948 2488 6160
<< metal4 >>
rect 285 9775 1485 10036
rect 2570 9770 3770 10036
rect 285 6171 1485 6273
rect 2769 6216 6781 6936
rect 1685 6171 2501 6173
rect 285 6160 2501 6171
rect 285 5948 2090 6160
rect 2488 5948 2501 6160
rect 285 4660 2501 5948
rect 6061 5601 6781 6216
use cc_via2_3cut  cc_via2_3cut_0
timestamp 1717772055
transform 0 1 -639040 -1 0 518654
box 517199 639873 517310 640172
use cc_via2_3cut  cc_via2_3cut_1
timestamp 1717772055
transform 0 1 -639448 -1 0 519454
box 517199 639873 517310 640172
use comparator_bias  comparator_bias_0
timestamp 1717776168
transform -1 0 518254 0 1 -639855
box 507866 646042 518182 649916
use comparator_core  comparator_core_0
timestamp 1717782065
transform 1 0 -506140 0 1 -641069
box 506214 638825 517124 647001
<< labels >>
flabel metal2 -140 1871 198 1971 0 FreeSans 1600 0 0 0 VINP
port 1 nsew
flabel metal2 -140 1636 198 1736 0 FreeSans 1600 0 0 0 VINM
port 0 nsew
flabel metal4 285 9775 1485 10036 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal4 2570 9770 3770 10036 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal2 11113 4077 11336 5865 0 FreeSans 1600 270 0 0 DVSS
port 6 nsew
flabel metal2 10902 3417 11337 3922 0 FreeSans 1600 0 0 0 DVDD
port 5 nsew
flabel metal2 10911 1738 11337 1838 0 FreeSans 1200 0 0 0 VOUT
port 7 nsew
<< end >>
