magic
tech sky130A
magscale 1 2
timestamp 1717725805
<< nmos >>
rect -1616 -531 -1016 469
rect -958 -531 -358 469
rect -300 -531 300 469
rect 358 -531 958 469
rect 1016 -531 1616 469
<< ndiff >>
rect -1674 457 -1616 469
rect -1674 -519 -1662 457
rect -1628 -519 -1616 457
rect -1674 -531 -1616 -519
rect -1016 457 -958 469
rect -1016 -519 -1004 457
rect -970 -519 -958 457
rect -1016 -531 -958 -519
rect -358 457 -300 469
rect -358 -519 -346 457
rect -312 -519 -300 457
rect -358 -531 -300 -519
rect 300 457 358 469
rect 300 -519 312 457
rect 346 -519 358 457
rect 300 -531 358 -519
rect 958 457 1016 469
rect 958 -519 970 457
rect 1004 -519 1016 457
rect 958 -531 1016 -519
rect 1616 457 1674 469
rect 1616 -519 1628 457
rect 1662 -519 1674 457
rect 1616 -531 1674 -519
<< ndiffc >>
rect -1662 -519 -1628 457
rect -1004 -519 -970 457
rect -346 -519 -312 457
rect 312 -519 346 457
rect 970 -519 1004 457
rect 1628 -519 1662 457
<< poly >>
rect -1616 541 -1016 557
rect -1616 507 -1600 541
rect -1032 507 -1016 541
rect -1616 469 -1016 507
rect -958 541 -358 557
rect -958 507 -942 541
rect -374 507 -358 541
rect -958 469 -358 507
rect -300 541 300 557
rect -300 507 -284 541
rect 284 507 300 541
rect -300 469 300 507
rect 358 541 958 557
rect 358 507 374 541
rect 942 507 958 541
rect 358 469 958 507
rect 1016 541 1616 557
rect 1016 507 1032 541
rect 1600 507 1616 541
rect 1016 469 1616 507
rect -1616 -557 -1016 -531
rect -958 -557 -358 -531
rect -300 -557 300 -531
rect 358 -557 958 -531
rect 1016 -557 1616 -531
<< polycont >>
rect -1600 507 -1032 541
rect -942 507 -374 541
rect -284 507 284 541
rect 374 507 942 541
rect 1032 507 1600 541
<< locali >>
rect -1616 507 -1600 541
rect -1032 507 -1016 541
rect -958 507 -942 541
rect -374 507 -358 541
rect -300 507 -284 541
rect 284 507 300 541
rect 358 507 374 541
rect 942 507 958 541
rect 1016 507 1032 541
rect 1600 507 1616 541
rect -1662 457 -1628 473
rect -1662 -535 -1628 -519
rect -1004 457 -970 473
rect -1004 -535 -970 -519
rect -346 457 -312 473
rect -346 -535 -312 -519
rect 312 457 346 473
rect 312 -535 346 -519
rect 970 457 1004 473
rect 970 -535 1004 -519
rect 1628 457 1662 473
rect 1628 -535 1662 -519
<< viali >>
rect -1600 507 -1032 541
rect -942 507 -374 541
rect -284 507 284 541
rect 374 507 942 541
rect 1032 507 1600 541
rect -1662 -519 -1628 457
rect -1004 -519 -970 457
rect -346 -519 -312 457
rect 312 -519 346 457
rect 970 -519 1004 457
rect 1628 -519 1662 457
<< metal1 >>
rect -1612 541 -1020 547
rect -1612 507 -1600 541
rect -1032 507 -1020 541
rect -1612 501 -1020 507
rect -954 541 -362 547
rect -954 507 -942 541
rect -374 507 -362 541
rect -954 501 -362 507
rect -296 541 296 547
rect -296 507 -284 541
rect 284 507 296 541
rect -296 501 296 507
rect 362 541 954 547
rect 362 507 374 541
rect 942 507 954 541
rect 362 501 954 507
rect 1020 541 1612 547
rect 1020 507 1032 541
rect 1600 507 1612 541
rect 1020 501 1612 507
rect -1668 457 -1622 469
rect -1668 -519 -1662 457
rect -1628 -519 -1622 457
rect -1668 -531 -1622 -519
rect -1010 457 -964 469
rect -1010 -519 -1004 457
rect -970 -519 -964 457
rect -1010 -531 -964 -519
rect -352 457 -306 469
rect -352 -519 -346 457
rect -312 -519 -306 457
rect -352 -531 -306 -519
rect 306 457 352 469
rect 306 -519 312 457
rect 346 -519 352 457
rect 306 -531 352 -519
rect 964 457 1010 469
rect 964 -519 970 457
rect 1004 -519 1010 457
rect 964 -531 1010 -519
rect 1622 457 1668 469
rect 1622 -519 1628 457
rect 1662 -519 1668 457
rect 1622 -531 1668 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 3 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
