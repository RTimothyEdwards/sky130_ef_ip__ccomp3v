magic
tech sky130A
magscale 1 2
timestamp 1717769754
<< checkpaint >>
rect 505457 643533 505524 643985
<< metal1 >>
rect 505457 643978 505524 643985
rect 505457 643533 505524 643540
<< via1 >>
rect 505457 643540 505524 643978
<< metal2 >>
rect 505457 643978 505524 643985
rect 505457 643533 505524 643540
<< end >>
