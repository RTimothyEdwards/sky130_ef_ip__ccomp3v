magic
tech sky130A
magscale 1 2
timestamp 1717772055
<< checkpaint >>
rect 517199 639873 517310 640172
<< metal2 >>
rect 517204 640160 517305 640172
rect 517204 639873 517305 639884
<< via2 >>
rect 517204 639884 517305 640160
<< metal3 >>
rect 517199 640160 517310 640172
rect 517199 639884 517204 640160
rect 517305 639884 517310 640160
rect 517199 639873 517310 639884
<< end >>
