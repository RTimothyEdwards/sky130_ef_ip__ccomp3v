magic
tech sky130A
magscale 1 2
timestamp 1717769384
<< checkpaint >>
rect 505947 645698 506014 646618
<< metal1 >>
rect 505947 646611 506014 646618
rect 505947 645698 506014 645705
<< via1 >>
rect 505947 645705 506014 646611
<< metal2 >>
rect 505947 646611 506014 646618
rect 505947 645698 506014 645705
<< end >>
