magic
tech sky130A
magscale 1 2
timestamp 1717725805
<< mvnmos >>
rect -1345 -531 -945 469
rect -887 -531 -487 469
rect -429 -531 -29 469
rect 29 -531 429 469
rect 487 -531 887 469
rect 945 -531 1345 469
<< mvndiff >>
rect -1403 457 -1345 469
rect -1403 -519 -1391 457
rect -1357 -519 -1345 457
rect -1403 -531 -1345 -519
rect -945 457 -887 469
rect -945 -519 -933 457
rect -899 -519 -887 457
rect -945 -531 -887 -519
rect -487 457 -429 469
rect -487 -519 -475 457
rect -441 -519 -429 457
rect -487 -531 -429 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 429 457 487 469
rect 429 -519 441 457
rect 475 -519 487 457
rect 429 -531 487 -519
rect 887 457 945 469
rect 887 -519 899 457
rect 933 -519 945 457
rect 887 -531 945 -519
rect 1345 457 1403 469
rect 1345 -519 1357 457
rect 1391 -519 1403 457
rect 1345 -531 1403 -519
<< mvndiffc >>
rect -1391 -519 -1357 457
rect -933 -519 -899 457
rect -475 -519 -441 457
rect -17 -519 17 457
rect 441 -519 475 457
rect 899 -519 933 457
rect 1357 -519 1391 457
<< poly >>
rect -1345 541 -945 557
rect -1345 507 -1329 541
rect -961 507 -945 541
rect -1345 469 -945 507
rect -887 541 -487 557
rect -887 507 -871 541
rect -503 507 -487 541
rect -887 469 -487 507
rect -429 541 -29 557
rect -429 507 -413 541
rect -45 507 -29 541
rect -429 469 -29 507
rect 29 541 429 557
rect 29 507 45 541
rect 413 507 429 541
rect 29 469 429 507
rect 487 541 887 557
rect 487 507 503 541
rect 871 507 887 541
rect 487 469 887 507
rect 945 541 1345 557
rect 945 507 961 541
rect 1329 507 1345 541
rect 945 469 1345 507
rect -1345 -557 -945 -531
rect -887 -557 -487 -531
rect -429 -557 -29 -531
rect 29 -557 429 -531
rect 487 -557 887 -531
rect 945 -557 1345 -531
<< polycont >>
rect -1329 507 -961 541
rect -871 507 -503 541
rect -413 507 -45 541
rect 45 507 413 541
rect 503 507 871 541
rect 961 507 1329 541
<< locali >>
rect -1345 507 -1329 541
rect -961 507 -945 541
rect -887 507 -871 541
rect -503 507 -487 541
rect -429 507 -413 541
rect -45 507 -29 541
rect 29 507 45 541
rect 413 507 429 541
rect 487 507 503 541
rect 871 507 887 541
rect 945 507 961 541
rect 1329 507 1345 541
rect -1391 457 -1357 473
rect -1391 -535 -1357 -519
rect -933 457 -899 473
rect -933 -535 -899 -519
rect -475 457 -441 473
rect -475 -535 -441 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 441 457 475 473
rect 441 -535 475 -519
rect 899 457 933 473
rect 899 -535 933 -519
rect 1357 457 1391 473
rect 1357 -535 1391 -519
<< viali >>
rect -1329 507 -961 541
rect -871 507 -503 541
rect -413 507 -45 541
rect 45 507 413 541
rect 503 507 871 541
rect 961 507 1329 541
rect -1391 -519 -1357 457
rect -933 -519 -899 457
rect -475 -519 -441 457
rect -17 -519 17 457
rect 441 -519 475 457
rect 899 -519 933 457
rect 1357 -519 1391 457
<< metal1 >>
rect -1341 541 -949 547
rect -1341 507 -1329 541
rect -961 507 -949 541
rect -1341 501 -949 507
rect -883 541 -491 547
rect -883 507 -871 541
rect -503 507 -491 541
rect -883 501 -491 507
rect -425 541 -33 547
rect -425 507 -413 541
rect -45 507 -33 541
rect -425 501 -33 507
rect 33 541 425 547
rect 33 507 45 541
rect 413 507 425 541
rect 33 501 425 507
rect 491 541 883 547
rect 491 507 503 541
rect 871 507 883 541
rect 491 501 883 507
rect 949 541 1341 547
rect 949 507 961 541
rect 1329 507 1341 541
rect 949 501 1341 507
rect -1397 457 -1351 469
rect -1397 -519 -1391 457
rect -1357 -519 -1351 457
rect -1397 -531 -1351 -519
rect -939 457 -893 469
rect -939 -519 -933 457
rect -899 -519 -893 457
rect -939 -531 -893 -519
rect -481 457 -435 469
rect -481 -519 -475 457
rect -441 -519 -435 457
rect -481 -531 -435 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 435 457 481 469
rect 435 -519 441 457
rect 475 -519 481 457
rect 435 -531 481 -519
rect 893 457 939 469
rect 893 -519 899 457
rect 933 -519 939 457
rect 893 -531 939 -519
rect 1351 457 1397 469
rect 1351 -519 1357 457
rect 1391 -519 1397 457
rect 1351 -531 1397 -519
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 2 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
