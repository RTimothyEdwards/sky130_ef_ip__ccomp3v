magic
tech sky130A
magscale 1 2
timestamp 1717765643
<< mvnmos >>
rect -1945 -531 -1345 469
rect -1287 -531 -687 469
rect -629 -531 -29 469
rect 29 -531 629 469
rect 687 -531 1287 469
rect 1345 -531 1945 469
<< mvndiff >>
rect -2003 457 -1945 469
rect -2003 -519 -1991 457
rect -1957 -519 -1945 457
rect -2003 -531 -1945 -519
rect -1345 457 -1287 469
rect -1345 -519 -1333 457
rect -1299 -519 -1287 457
rect -1345 -531 -1287 -519
rect -687 457 -629 469
rect -687 -519 -675 457
rect -641 -519 -629 457
rect -687 -531 -629 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 629 457 687 469
rect 629 -519 641 457
rect 675 -519 687 457
rect 629 -531 687 -519
rect 1287 457 1345 469
rect 1287 -519 1299 457
rect 1333 -519 1345 457
rect 1287 -531 1345 -519
rect 1945 457 2003 469
rect 1945 -519 1957 457
rect 1991 -519 2003 457
rect 1945 -531 2003 -519
<< mvndiffc >>
rect -1991 -519 -1957 457
rect -1333 -519 -1299 457
rect -675 -519 -641 457
rect -17 -519 17 457
rect 641 -519 675 457
rect 1299 -519 1333 457
rect 1957 -519 1991 457
<< poly >>
rect -1945 541 -1345 557
rect -1945 507 -1929 541
rect -1361 507 -1345 541
rect -1945 469 -1345 507
rect -1287 541 -687 557
rect -1287 507 -1271 541
rect -703 507 -687 541
rect -1287 469 -687 507
rect -629 541 -29 557
rect -629 507 -613 541
rect -45 507 -29 541
rect -629 469 -29 507
rect 29 541 629 557
rect 29 507 45 541
rect 613 507 629 541
rect 29 469 629 507
rect 687 541 1287 557
rect 687 507 703 541
rect 1271 507 1287 541
rect 687 469 1287 507
rect 1345 541 1945 557
rect 1345 507 1361 541
rect 1929 507 1945 541
rect 1345 469 1945 507
rect -1945 -557 -1345 -531
rect -1287 -557 -687 -531
rect -629 -557 -29 -531
rect 29 -557 629 -531
rect 687 -557 1287 -531
rect 1345 -557 1945 -531
<< polycont >>
rect -1929 507 -1361 541
rect -1271 507 -703 541
rect -613 507 -45 541
rect 45 507 613 541
rect 703 507 1271 541
rect 1361 507 1929 541
<< locali >>
rect -1945 507 -1929 541
rect -1361 507 -1345 541
rect -1287 507 -1271 541
rect -703 507 -687 541
rect -629 507 -613 541
rect -45 507 -29 541
rect 29 507 45 541
rect 613 507 629 541
rect 687 507 703 541
rect 1271 507 1287 541
rect 1345 507 1361 541
rect 1929 507 1945 541
rect -1991 457 -1957 473
rect -1991 -535 -1957 -519
rect -1333 457 -1299 473
rect -1333 -535 -1299 -519
rect -675 457 -641 473
rect -675 -535 -641 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 641 457 675 473
rect 641 -535 675 -519
rect 1299 457 1333 473
rect 1299 -535 1333 -519
rect 1957 457 1991 473
rect 1957 -535 1991 -519
<< viali >>
rect -1929 507 -1361 541
rect -1271 507 -703 541
rect -613 507 -45 541
rect 45 507 613 541
rect 703 507 1271 541
rect 1361 507 1929 541
rect -1991 -519 -1957 457
rect -1333 -519 -1299 457
rect -675 -519 -641 457
rect -17 -519 17 457
rect 641 -519 675 457
rect 1299 -519 1333 457
rect 1957 -519 1991 457
<< metal1 >>
rect -1941 541 -1349 547
rect -1941 507 -1929 541
rect -1361 507 -1349 541
rect -1941 501 -1349 507
rect -1283 541 -691 547
rect -1283 507 -1271 541
rect -703 507 -691 541
rect -1283 501 -691 507
rect -625 541 -33 547
rect -625 507 -613 541
rect -45 507 -33 541
rect -625 501 -33 507
rect 33 541 625 547
rect 33 507 45 541
rect 613 507 625 541
rect 33 501 625 507
rect 691 541 1283 547
rect 691 507 703 541
rect 1271 507 1283 541
rect 691 501 1283 507
rect 1349 541 1941 547
rect 1349 507 1361 541
rect 1929 507 1941 541
rect 1349 501 1941 507
rect -1997 457 -1951 469
rect -1997 -519 -1991 457
rect -1957 -519 -1951 457
rect -1997 -531 -1951 -519
rect -1339 457 -1293 469
rect -1339 -519 -1333 457
rect -1299 -519 -1293 457
rect -1339 -531 -1293 -519
rect -681 457 -635 469
rect -681 -519 -675 457
rect -641 -519 -635 457
rect -681 -531 -635 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 635 457 681 469
rect 635 -519 641 457
rect 675 -519 681 457
rect 635 -531 681 -519
rect 1293 457 1339 469
rect 1293 -519 1299 457
rect 1333 -519 1339 457
rect 1293 -531 1339 -519
rect 1951 457 1997 469
rect 1951 -519 1957 457
rect 1991 -519 1997 457
rect 1951 -531 1997 -519
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 3 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
