magic
tech sky130A
magscale 1 2
timestamp 1717725805
<< nwell >>
rect -1439 -564 1439 598
<< pmos >>
rect -1345 -464 -945 536
rect -887 -464 -487 536
rect -429 -464 -29 536
rect 29 -464 429 536
rect 487 -464 887 536
rect 945 -464 1345 536
<< pdiff >>
rect -1403 524 -1345 536
rect -1403 -452 -1391 524
rect -1357 -452 -1345 524
rect -1403 -464 -1345 -452
rect -945 524 -887 536
rect -945 -452 -933 524
rect -899 -452 -887 524
rect -945 -464 -887 -452
rect -487 524 -429 536
rect -487 -452 -475 524
rect -441 -452 -429 524
rect -487 -464 -429 -452
rect -29 524 29 536
rect -29 -452 -17 524
rect 17 -452 29 524
rect -29 -464 29 -452
rect 429 524 487 536
rect 429 -452 441 524
rect 475 -452 487 524
rect 429 -464 487 -452
rect 887 524 945 536
rect 887 -452 899 524
rect 933 -452 945 524
rect 887 -464 945 -452
rect 1345 524 1403 536
rect 1345 -452 1357 524
rect 1391 -452 1403 524
rect 1345 -464 1403 -452
<< pdiffc >>
rect -1391 -452 -1357 524
rect -933 -452 -899 524
rect -475 -452 -441 524
rect -17 -452 17 524
rect 441 -452 475 524
rect 899 -452 933 524
rect 1357 -452 1391 524
<< poly >>
rect -1345 536 -945 562
rect -887 536 -487 562
rect -429 536 -29 562
rect 29 536 429 562
rect 487 536 887 562
rect 945 536 1345 562
rect -1345 -511 -945 -464
rect -1345 -545 -1329 -511
rect -961 -545 -945 -511
rect -1345 -561 -945 -545
rect -887 -511 -487 -464
rect -887 -545 -871 -511
rect -503 -545 -487 -511
rect -887 -561 -487 -545
rect -429 -511 -29 -464
rect -429 -545 -413 -511
rect -45 -545 -29 -511
rect -429 -561 -29 -545
rect 29 -511 429 -464
rect 29 -545 45 -511
rect 413 -545 429 -511
rect 29 -561 429 -545
rect 487 -511 887 -464
rect 487 -545 503 -511
rect 871 -545 887 -511
rect 487 -561 887 -545
rect 945 -511 1345 -464
rect 945 -545 961 -511
rect 1329 -545 1345 -511
rect 945 -561 1345 -545
<< polycont >>
rect -1329 -545 -961 -511
rect -871 -545 -503 -511
rect -413 -545 -45 -511
rect 45 -545 413 -511
rect 503 -545 871 -511
rect 961 -545 1329 -511
<< locali >>
rect -1391 524 -1357 540
rect -1391 -468 -1357 -452
rect -933 524 -899 540
rect -933 -468 -899 -452
rect -475 524 -441 540
rect -475 -468 -441 -452
rect -17 524 17 540
rect -17 -468 17 -452
rect 441 524 475 540
rect 441 -468 475 -452
rect 899 524 933 540
rect 899 -468 933 -452
rect 1357 524 1391 540
rect 1357 -468 1391 -452
rect -1345 -545 -1329 -511
rect -961 -545 -945 -511
rect -887 -545 -871 -511
rect -503 -545 -487 -511
rect -429 -545 -413 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 413 -545 429 -511
rect 487 -545 503 -511
rect 871 -545 887 -511
rect 945 -545 961 -511
rect 1329 -545 1345 -511
<< viali >>
rect -1391 -452 -1357 524
rect -933 -452 -899 524
rect -475 -452 -441 524
rect -17 -452 17 524
rect 441 -452 475 524
rect 899 -452 933 524
rect 1357 -452 1391 524
rect -1329 -545 -961 -511
rect -871 -545 -503 -511
rect -413 -545 -45 -511
rect 45 -545 413 -511
rect 503 -545 871 -511
rect 961 -545 1329 -511
<< metal1 >>
rect -1397 524 -1351 536
rect -1397 -452 -1391 524
rect -1357 -452 -1351 524
rect -1397 -464 -1351 -452
rect -939 524 -893 536
rect -939 -452 -933 524
rect -899 -452 -893 524
rect -939 -464 -893 -452
rect -481 524 -435 536
rect -481 -452 -475 524
rect -441 -452 -435 524
rect -481 -464 -435 -452
rect -23 524 23 536
rect -23 -452 -17 524
rect 17 -452 23 524
rect -23 -464 23 -452
rect 435 524 481 536
rect 435 -452 441 524
rect 475 -452 481 524
rect 435 -464 481 -452
rect 893 524 939 536
rect 893 -452 899 524
rect 933 -452 939 524
rect 893 -464 939 -452
rect 1351 524 1397 536
rect 1351 -452 1357 524
rect 1391 -452 1397 524
rect 1351 -464 1397 -452
rect -1341 -511 -949 -505
rect -1341 -545 -1329 -511
rect -961 -545 -949 -511
rect -1341 -551 -949 -545
rect -883 -511 -491 -505
rect -883 -545 -871 -511
rect -503 -545 -491 -511
rect -883 -551 -491 -545
rect -425 -511 -33 -505
rect -425 -545 -413 -511
rect -45 -545 -33 -511
rect -425 -551 -33 -545
rect 33 -511 425 -505
rect 33 -545 45 -511
rect 413 -545 425 -511
rect 33 -551 425 -545
rect 491 -511 883 -505
rect 491 -545 503 -511
rect 871 -545 883 -511
rect 491 -551 883 -545
rect 949 -511 1341 -505
rect 949 -545 961 -511
rect 1329 -545 1341 -511
rect 949 -551 1341 -545
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 2 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
