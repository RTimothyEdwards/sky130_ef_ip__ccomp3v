magic
tech sky130A
magscale 1 2
timestamp 1731000523
<< pwell >>
rect -428 -1327 428 1327
<< mvnmos >>
rect -200 109 200 1069
rect -200 -1069 200 -109
<< mvndiff >>
rect -258 1057 -200 1069
rect -258 121 -246 1057
rect -212 121 -200 1057
rect -258 109 -200 121
rect 200 1057 258 1069
rect 200 121 212 1057
rect 246 121 258 1057
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -1057 -246 -121
rect -212 -1057 -200 -121
rect -258 -1069 -200 -1057
rect 200 -121 258 -109
rect 200 -1057 212 -121
rect 246 -1057 258 -121
rect 200 -1069 258 -1057
<< mvndiffc >>
rect -246 121 -212 1057
rect 212 121 246 1057
rect -246 -1057 -212 -121
rect 212 -1057 246 -121
<< mvpsubdiff >>
rect -392 1279 392 1291
rect -392 1245 -284 1279
rect 284 1245 392 1279
rect -392 1233 392 1245
rect -392 1183 -334 1233
rect -392 -1183 -380 1183
rect -346 -1183 -334 1183
rect 334 1183 392 1233
rect -392 -1233 -334 -1183
rect 334 -1183 346 1183
rect 380 -1183 392 1183
rect 334 -1233 392 -1183
rect -392 -1245 392 -1233
rect -392 -1279 -284 -1245
rect 284 -1279 392 -1245
rect -392 -1291 392 -1279
<< mvpsubdiffcont >>
rect -284 1245 284 1279
rect -380 -1183 -346 1183
rect 346 -1183 380 1183
rect -284 -1279 284 -1245
<< poly >>
rect -200 1141 200 1157
rect -200 1107 -184 1141
rect 184 1107 200 1141
rect -200 1069 200 1107
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -1107 200 -1069
rect -200 -1141 -184 -1107
rect 184 -1141 200 -1107
rect -200 -1157 200 -1141
<< polycont >>
rect -184 1107 184 1141
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -1141 184 -1107
<< locali >>
rect -380 1245 -284 1279
rect 284 1245 380 1279
rect -380 1183 -346 1245
rect 346 1183 380 1245
rect -200 1107 -184 1141
rect 184 1107 200 1141
rect -246 1057 -212 1073
rect -246 105 -212 121
rect 212 1057 246 1073
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -1073 -212 -1057
rect 212 -121 246 -105
rect 212 -1073 246 -1057
rect -200 -1141 -184 -1107
rect 184 -1141 200 -1107
rect -380 -1245 -346 -1183
rect 346 -1245 380 -1183
rect -380 -1279 -284 -1245
rect 284 -1279 380 -1245
<< viali >>
rect -184 1107 184 1141
rect -246 121 -212 1057
rect 212 121 246 1057
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -1057 -212 -121
rect 212 -1057 246 -121
rect -184 -1141 184 -1107
<< metal1 >>
rect -196 1141 196 1147
rect -196 1107 -184 1141
rect 184 1107 196 1141
rect -196 1101 196 1107
rect -252 1057 -206 1069
rect -252 121 -246 1057
rect -212 121 -206 1057
rect -252 109 -206 121
rect 206 1057 252 1069
rect 206 121 212 1057
rect 246 121 252 1057
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -1057 -246 -121
rect -212 -1057 -206 -121
rect -252 -1069 -206 -1057
rect 206 -121 252 -109
rect 206 -1057 212 -121
rect 246 -1057 252 -121
rect 206 -1069 252 -1057
rect -196 -1107 196 -1101
rect -196 -1141 -184 -1107
rect 184 -1141 196 -1107
rect -196 -1147 196 -1141
<< properties >>
string FIXED_BBOX -363 -1262 363 1262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.8 l 2.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
