magic
tech sky130A
magscale 1 2
timestamp 1731000523
<< pwell >>
rect -428 -1367 428 1367
<< mvnmos >>
rect -200 109 200 1109
rect -200 -1109 200 -109
<< mvndiff >>
rect -258 1097 -200 1109
rect -258 121 -246 1097
rect -212 121 -200 1097
rect -258 109 -200 121
rect 200 1097 258 1109
rect 200 121 212 1097
rect 246 121 258 1097
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -1097 -246 -121
rect -212 -1097 -200 -121
rect -258 -1109 -200 -1097
rect 200 -121 258 -109
rect 200 -1097 212 -121
rect 246 -1097 258 -121
rect 200 -1109 258 -1097
<< mvndiffc >>
rect -246 121 -212 1097
rect 212 121 246 1097
rect -246 -1097 -212 -121
rect 212 -1097 246 -121
<< mvpsubdiff >>
rect -392 1319 392 1331
rect -392 1285 -284 1319
rect 284 1285 392 1319
rect -392 1273 392 1285
rect -392 1223 -334 1273
rect -392 -1223 -380 1223
rect -346 -1223 -334 1223
rect 334 1223 392 1273
rect -392 -1273 -334 -1223
rect 334 -1223 346 1223
rect 380 -1223 392 1223
rect 334 -1273 392 -1223
rect -392 -1285 392 -1273
rect -392 -1319 -284 -1285
rect 284 -1319 392 -1285
rect -392 -1331 392 -1319
<< mvpsubdiffcont >>
rect -284 1285 284 1319
rect -380 -1223 -346 1223
rect 346 -1223 380 1223
rect -284 -1319 284 -1285
<< poly >>
rect -200 1181 200 1197
rect -200 1147 -184 1181
rect 184 1147 200 1181
rect -200 1109 200 1147
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -1147 200 -1109
rect -200 -1181 -184 -1147
rect 184 -1181 200 -1147
rect -200 -1197 200 -1181
<< polycont >>
rect -184 1147 184 1181
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -1181 184 -1147
<< locali >>
rect -380 1285 -284 1319
rect 284 1285 380 1319
rect -380 1223 -346 1285
rect 346 1223 380 1285
rect -200 1147 -184 1181
rect 184 1147 200 1181
rect -246 1097 -212 1113
rect -246 105 -212 121
rect 212 1097 246 1113
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -1113 -212 -1097
rect 212 -121 246 -105
rect 212 -1113 246 -1097
rect -200 -1181 -184 -1147
rect 184 -1181 200 -1147
rect -380 -1285 -346 -1223
rect 346 -1285 380 -1223
rect -380 -1319 -284 -1285
rect 284 -1319 380 -1285
<< viali >>
rect -184 1147 184 1181
rect -246 121 -212 1097
rect 212 121 246 1097
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -1097 -212 -121
rect 212 -1097 246 -121
rect -184 -1181 184 -1147
<< metal1 >>
rect -196 1181 196 1187
rect -196 1147 -184 1181
rect 184 1147 196 1181
rect -196 1141 196 1147
rect -252 1097 -206 1109
rect -252 121 -246 1097
rect -212 121 -206 1097
rect -252 109 -206 121
rect 206 1097 252 1109
rect 206 121 212 1097
rect 246 121 252 1097
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -1097 -246 -121
rect -212 -1097 -206 -121
rect -252 -1109 -206 -1097
rect 206 -121 252 -109
rect 206 -1097 212 -121
rect 246 -1097 252 -121
rect 206 -1109 252 -1097
rect -196 -1147 196 -1141
rect -196 -1181 -184 -1147
rect 184 -1181 196 -1147
rect -196 -1187 196 -1181
<< properties >>
string FIXED_BBOX -363 -1302 363 1302
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 2.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
