magic
tech sky130A
magscale 1 2
timestamp 1731000523
<< pwell >>
rect -328 -6239 328 6239
<< mvnnmos >>
rect -100 4981 100 5981
rect -100 3763 100 4763
rect -100 2545 100 3545
rect -100 1327 100 2327
rect -100 109 100 1109
rect -100 -1109 100 -109
rect -100 -2327 100 -1327
rect -100 -3545 100 -2545
rect -100 -4763 100 -3763
rect -100 -5981 100 -4981
<< mvndiff >>
rect -158 5969 -100 5981
rect -158 4993 -146 5969
rect -112 4993 -100 5969
rect -158 4981 -100 4993
rect 100 5969 158 5981
rect 100 4993 112 5969
rect 146 4993 158 5969
rect 100 4981 158 4993
rect -158 4751 -100 4763
rect -158 3775 -146 4751
rect -112 3775 -100 4751
rect -158 3763 -100 3775
rect 100 4751 158 4763
rect 100 3775 112 4751
rect 146 3775 158 4751
rect 100 3763 158 3775
rect -158 3533 -100 3545
rect -158 2557 -146 3533
rect -112 2557 -100 3533
rect -158 2545 -100 2557
rect 100 3533 158 3545
rect 100 2557 112 3533
rect 146 2557 158 3533
rect 100 2545 158 2557
rect -158 2315 -100 2327
rect -158 1339 -146 2315
rect -112 1339 -100 2315
rect -158 1327 -100 1339
rect 100 2315 158 2327
rect 100 1339 112 2315
rect 146 1339 158 2315
rect 100 1327 158 1339
rect -158 1097 -100 1109
rect -158 121 -146 1097
rect -112 121 -100 1097
rect -158 109 -100 121
rect 100 1097 158 1109
rect 100 121 112 1097
rect 146 121 158 1097
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1097 -146 -121
rect -112 -1097 -100 -121
rect -158 -1109 -100 -1097
rect 100 -121 158 -109
rect 100 -1097 112 -121
rect 146 -1097 158 -121
rect 100 -1109 158 -1097
rect -158 -1339 -100 -1327
rect -158 -2315 -146 -1339
rect -112 -2315 -100 -1339
rect -158 -2327 -100 -2315
rect 100 -1339 158 -1327
rect 100 -2315 112 -1339
rect 146 -2315 158 -1339
rect 100 -2327 158 -2315
rect -158 -2557 -100 -2545
rect -158 -3533 -146 -2557
rect -112 -3533 -100 -2557
rect -158 -3545 -100 -3533
rect 100 -2557 158 -2545
rect 100 -3533 112 -2557
rect 146 -3533 158 -2557
rect 100 -3545 158 -3533
rect -158 -3775 -100 -3763
rect -158 -4751 -146 -3775
rect -112 -4751 -100 -3775
rect -158 -4763 -100 -4751
rect 100 -3775 158 -3763
rect 100 -4751 112 -3775
rect 146 -4751 158 -3775
rect 100 -4763 158 -4751
rect -158 -4993 -100 -4981
rect -158 -5969 -146 -4993
rect -112 -5969 -100 -4993
rect -158 -5981 -100 -5969
rect 100 -4993 158 -4981
rect 100 -5969 112 -4993
rect 146 -5969 158 -4993
rect 100 -5981 158 -5969
<< mvndiffc >>
rect -146 4993 -112 5969
rect 112 4993 146 5969
rect -146 3775 -112 4751
rect 112 3775 146 4751
rect -146 2557 -112 3533
rect 112 2557 146 3533
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect -146 121 -112 1097
rect 112 121 146 1097
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect -146 -3533 -112 -2557
rect 112 -3533 146 -2557
rect -146 -4751 -112 -3775
rect 112 -4751 146 -3775
rect -146 -5969 -112 -4993
rect 112 -5969 146 -4993
<< mvpsubdiff >>
rect -292 6191 292 6203
rect -292 6157 -184 6191
rect 184 6157 292 6191
rect -292 6145 292 6157
rect -292 6095 -234 6145
rect -292 -6095 -280 6095
rect -246 -6095 -234 6095
rect 234 6095 292 6145
rect -292 -6145 -234 -6095
rect 234 -6095 246 6095
rect 280 -6095 292 6095
rect 234 -6145 292 -6095
rect -292 -6157 292 -6145
rect -292 -6191 -184 -6157
rect 184 -6191 292 -6157
rect -292 -6203 292 -6191
<< mvpsubdiffcont >>
rect -184 6157 184 6191
rect -280 -6095 -246 6095
rect 246 -6095 280 6095
rect -184 -6191 184 -6157
<< poly >>
rect -100 6053 100 6069
rect -100 6019 -84 6053
rect 84 6019 100 6053
rect -100 5981 100 6019
rect -100 4943 100 4981
rect -100 4909 -84 4943
rect 84 4909 100 4943
rect -100 4893 100 4909
rect -100 4835 100 4851
rect -100 4801 -84 4835
rect 84 4801 100 4835
rect -100 4763 100 4801
rect -100 3725 100 3763
rect -100 3691 -84 3725
rect 84 3691 100 3725
rect -100 3675 100 3691
rect -100 3617 100 3633
rect -100 3583 -84 3617
rect 84 3583 100 3617
rect -100 3545 100 3583
rect -100 2507 100 2545
rect -100 2473 -84 2507
rect 84 2473 100 2507
rect -100 2457 100 2473
rect -100 2399 100 2415
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -100 2327 100 2365
rect -100 1289 100 1327
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1239 100 1255
rect -100 1181 100 1197
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -100 1109 100 1147
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1147 100 -1109
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1197 100 -1181
rect -100 -1255 100 -1239
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -100 -1327 100 -1289
rect -100 -2365 100 -2327
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2415 100 -2399
rect -100 -2473 100 -2457
rect -100 -2507 -84 -2473
rect 84 -2507 100 -2473
rect -100 -2545 100 -2507
rect -100 -3583 100 -3545
rect -100 -3617 -84 -3583
rect 84 -3617 100 -3583
rect -100 -3633 100 -3617
rect -100 -3691 100 -3675
rect -100 -3725 -84 -3691
rect 84 -3725 100 -3691
rect -100 -3763 100 -3725
rect -100 -4801 100 -4763
rect -100 -4835 -84 -4801
rect 84 -4835 100 -4801
rect -100 -4851 100 -4835
rect -100 -4909 100 -4893
rect -100 -4943 -84 -4909
rect 84 -4943 100 -4909
rect -100 -4981 100 -4943
rect -100 -6019 100 -5981
rect -100 -6053 -84 -6019
rect 84 -6053 100 -6019
rect -100 -6069 100 -6053
<< polycont >>
rect -84 6019 84 6053
rect -84 4909 84 4943
rect -84 4801 84 4835
rect -84 3691 84 3725
rect -84 3583 84 3617
rect -84 2473 84 2507
rect -84 2365 84 2399
rect -84 1255 84 1289
rect -84 1147 84 1181
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1181 84 -1147
rect -84 -1289 84 -1255
rect -84 -2399 84 -2365
rect -84 -2507 84 -2473
rect -84 -3617 84 -3583
rect -84 -3725 84 -3691
rect -84 -4835 84 -4801
rect -84 -4943 84 -4909
rect -84 -6053 84 -6019
<< locali >>
rect -280 6157 -184 6191
rect 184 6157 280 6191
rect -280 6095 -246 6157
rect 246 6095 280 6157
rect -100 6019 -84 6053
rect 84 6019 100 6053
rect -146 5969 -112 5985
rect -146 4977 -112 4993
rect 112 5969 146 5985
rect 112 4977 146 4993
rect -100 4909 -84 4943
rect 84 4909 100 4943
rect -100 4801 -84 4835
rect 84 4801 100 4835
rect -146 4751 -112 4767
rect -146 3759 -112 3775
rect 112 4751 146 4767
rect 112 3759 146 3775
rect -100 3691 -84 3725
rect 84 3691 100 3725
rect -100 3583 -84 3617
rect 84 3583 100 3617
rect -146 3533 -112 3549
rect -146 2541 -112 2557
rect 112 3533 146 3549
rect 112 2541 146 2557
rect -100 2473 -84 2507
rect 84 2473 100 2507
rect -100 2365 -84 2399
rect 84 2365 100 2399
rect -146 2315 -112 2331
rect -146 1323 -112 1339
rect 112 2315 146 2331
rect 112 1323 146 1339
rect -100 1255 -84 1289
rect 84 1255 100 1289
rect -100 1147 -84 1181
rect 84 1147 100 1181
rect -146 1097 -112 1113
rect -146 105 -112 121
rect 112 1097 146 1113
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1113 -112 -1097
rect 112 -121 146 -105
rect 112 -1113 146 -1097
rect -100 -1181 -84 -1147
rect 84 -1181 100 -1147
rect -100 -1289 -84 -1255
rect 84 -1289 100 -1255
rect -146 -1339 -112 -1323
rect -146 -2331 -112 -2315
rect 112 -1339 146 -1323
rect 112 -2331 146 -2315
rect -100 -2399 -84 -2365
rect 84 -2399 100 -2365
rect -100 -2507 -84 -2473
rect 84 -2507 100 -2473
rect -146 -2557 -112 -2541
rect -146 -3549 -112 -3533
rect 112 -2557 146 -2541
rect 112 -3549 146 -3533
rect -100 -3617 -84 -3583
rect 84 -3617 100 -3583
rect -100 -3725 -84 -3691
rect 84 -3725 100 -3691
rect -146 -3775 -112 -3759
rect -146 -4767 -112 -4751
rect 112 -3775 146 -3759
rect 112 -4767 146 -4751
rect -100 -4835 -84 -4801
rect 84 -4835 100 -4801
rect -100 -4943 -84 -4909
rect 84 -4943 100 -4909
rect -146 -4993 -112 -4977
rect -146 -5985 -112 -5969
rect 112 -4993 146 -4977
rect 112 -5985 146 -5969
rect -100 -6053 -84 -6019
rect 84 -6053 100 -6019
rect -280 -6157 -246 -6095
rect 246 -6157 280 -6095
rect -280 -6191 -184 -6157
rect 184 -6191 280 -6157
<< viali >>
rect -84 6019 84 6053
rect -146 4993 -112 5969
rect 112 4993 146 5969
rect -84 4909 84 4943
rect -84 4801 84 4835
rect -146 3775 -112 4751
rect 112 3775 146 4751
rect -84 3691 84 3725
rect -84 3583 84 3617
rect -146 2557 -112 3533
rect 112 2557 146 3533
rect -84 2473 84 2507
rect -84 2365 84 2399
rect -146 1339 -112 2315
rect 112 1339 146 2315
rect -84 1255 84 1289
rect -84 1147 84 1181
rect -146 121 -112 1097
rect 112 121 146 1097
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1097 -112 -121
rect 112 -1097 146 -121
rect -84 -1181 84 -1147
rect -84 -1289 84 -1255
rect -146 -2315 -112 -1339
rect 112 -2315 146 -1339
rect -84 -2399 84 -2365
rect -84 -2507 84 -2473
rect -146 -3533 -112 -2557
rect 112 -3533 146 -2557
rect -84 -3617 84 -3583
rect -84 -3725 84 -3691
rect -146 -4751 -112 -3775
rect 112 -4751 146 -3775
rect -84 -4835 84 -4801
rect -84 -4943 84 -4909
rect -146 -5969 -112 -4993
rect 112 -5969 146 -4993
rect -84 -6053 84 -6019
<< metal1 >>
rect -96 6053 96 6059
rect -96 6019 -84 6053
rect 84 6019 96 6053
rect -96 6013 96 6019
rect -152 5969 -106 5981
rect -152 4993 -146 5969
rect -112 4993 -106 5969
rect -152 4981 -106 4993
rect 106 5969 152 5981
rect 106 4993 112 5969
rect 146 4993 152 5969
rect 106 4981 152 4993
rect -96 4943 96 4949
rect -96 4909 -84 4943
rect 84 4909 96 4943
rect -96 4903 96 4909
rect -96 4835 96 4841
rect -96 4801 -84 4835
rect 84 4801 96 4835
rect -96 4795 96 4801
rect -152 4751 -106 4763
rect -152 3775 -146 4751
rect -112 3775 -106 4751
rect -152 3763 -106 3775
rect 106 4751 152 4763
rect 106 3775 112 4751
rect 146 3775 152 4751
rect 106 3763 152 3775
rect -96 3725 96 3731
rect -96 3691 -84 3725
rect 84 3691 96 3725
rect -96 3685 96 3691
rect -96 3617 96 3623
rect -96 3583 -84 3617
rect 84 3583 96 3617
rect -96 3577 96 3583
rect -152 3533 -106 3545
rect -152 2557 -146 3533
rect -112 2557 -106 3533
rect -152 2545 -106 2557
rect 106 3533 152 3545
rect 106 2557 112 3533
rect 146 2557 152 3533
rect 106 2545 152 2557
rect -96 2507 96 2513
rect -96 2473 -84 2507
rect 84 2473 96 2507
rect -96 2467 96 2473
rect -96 2399 96 2405
rect -96 2365 -84 2399
rect 84 2365 96 2399
rect -96 2359 96 2365
rect -152 2315 -106 2327
rect -152 1339 -146 2315
rect -112 1339 -106 2315
rect -152 1327 -106 1339
rect 106 2315 152 2327
rect 106 1339 112 2315
rect 146 1339 152 2315
rect 106 1327 152 1339
rect -96 1289 96 1295
rect -96 1255 -84 1289
rect 84 1255 96 1289
rect -96 1249 96 1255
rect -96 1181 96 1187
rect -96 1147 -84 1181
rect 84 1147 96 1181
rect -96 1141 96 1147
rect -152 1097 -106 1109
rect -152 121 -146 1097
rect -112 121 -106 1097
rect -152 109 -106 121
rect 106 1097 152 1109
rect 106 121 112 1097
rect 146 121 152 1097
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -1097 -146 -121
rect -112 -1097 -106 -121
rect -152 -1109 -106 -1097
rect 106 -121 152 -109
rect 106 -1097 112 -121
rect 146 -1097 152 -121
rect 106 -1109 152 -1097
rect -96 -1147 96 -1141
rect -96 -1181 -84 -1147
rect 84 -1181 96 -1147
rect -96 -1187 96 -1181
rect -96 -1255 96 -1249
rect -96 -1289 -84 -1255
rect 84 -1289 96 -1255
rect -96 -1295 96 -1289
rect -152 -1339 -106 -1327
rect -152 -2315 -146 -1339
rect -112 -2315 -106 -1339
rect -152 -2327 -106 -2315
rect 106 -1339 152 -1327
rect 106 -2315 112 -1339
rect 146 -2315 152 -1339
rect 106 -2327 152 -2315
rect -96 -2365 96 -2359
rect -96 -2399 -84 -2365
rect 84 -2399 96 -2365
rect -96 -2405 96 -2399
rect -96 -2473 96 -2467
rect -96 -2507 -84 -2473
rect 84 -2507 96 -2473
rect -96 -2513 96 -2507
rect -152 -2557 -106 -2545
rect -152 -3533 -146 -2557
rect -112 -3533 -106 -2557
rect -152 -3545 -106 -3533
rect 106 -2557 152 -2545
rect 106 -3533 112 -2557
rect 146 -3533 152 -2557
rect 106 -3545 152 -3533
rect -96 -3583 96 -3577
rect -96 -3617 -84 -3583
rect 84 -3617 96 -3583
rect -96 -3623 96 -3617
rect -96 -3691 96 -3685
rect -96 -3725 -84 -3691
rect 84 -3725 96 -3691
rect -96 -3731 96 -3725
rect -152 -3775 -106 -3763
rect -152 -4751 -146 -3775
rect -112 -4751 -106 -3775
rect -152 -4763 -106 -4751
rect 106 -3775 152 -3763
rect 106 -4751 112 -3775
rect 146 -4751 152 -3775
rect 106 -4763 152 -4751
rect -96 -4801 96 -4795
rect -96 -4835 -84 -4801
rect 84 -4835 96 -4801
rect -96 -4841 96 -4835
rect -96 -4909 96 -4903
rect -96 -4943 -84 -4909
rect 84 -4943 96 -4909
rect -96 -4949 96 -4943
rect -152 -4993 -106 -4981
rect -152 -5969 -146 -4993
rect -112 -5969 -106 -4993
rect -152 -5981 -106 -5969
rect 106 -4993 152 -4981
rect 106 -5969 112 -4993
rect 146 -5969 152 -4993
rect 106 -5981 152 -5969
rect -96 -6019 96 -6013
rect -96 -6053 -84 -6019
rect 84 -6053 96 -6019
rect -96 -6059 96 -6053
<< properties >>
string FIXED_BBOX -263 -6174 263 6174
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 5.0 l 1.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
