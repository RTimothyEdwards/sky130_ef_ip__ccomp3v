magic
tech sky130A
magscale 1 2
timestamp 1717725805
<< nmos >>
rect -379 -531 -29 469
rect 29 -531 379 469
<< ndiff >>
rect -437 457 -379 469
rect -437 -519 -425 457
rect -391 -519 -379 457
rect -437 -531 -379 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 379 457 437 469
rect 379 -519 391 457
rect 425 -519 437 457
rect 379 -531 437 -519
<< ndiffc >>
rect -425 -519 -391 457
rect -17 -519 17 457
rect 391 -519 425 457
<< poly >>
rect -379 541 -29 557
rect -379 507 -363 541
rect -45 507 -29 541
rect -379 469 -29 507
rect 29 541 379 557
rect 29 507 45 541
rect 363 507 379 541
rect 29 469 379 507
rect -379 -557 -29 -531
rect 29 -557 379 -531
<< polycont >>
rect -363 507 -45 541
rect 45 507 363 541
<< locali >>
rect -379 507 -363 541
rect -45 507 -29 541
rect 29 507 45 541
rect 363 507 379 541
rect -425 457 -391 473
rect -425 -535 -391 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 391 457 425 473
rect 391 -535 425 -519
<< viali >>
rect -363 507 -45 541
rect 45 507 363 541
rect -425 -519 -391 457
rect -17 -519 17 457
rect 391 -519 425 457
<< metal1 >>
rect -375 541 -33 547
rect -375 507 -363 541
rect -45 507 -33 541
rect -375 501 -33 507
rect 33 541 375 547
rect 33 507 45 541
rect 363 507 375 541
rect 33 501 375 507
rect -431 457 -385 469
rect -431 -519 -425 457
rect -391 -519 -385 457
rect -431 -531 -385 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 385 457 431 469
rect 385 -519 391 457
rect 425 -519 431 457
rect 385 -531 431 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1.75 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
