magic
tech sky130A
magscale 1 2
timestamp 1721179627
<< dnwell >>
rect -91 6072 10341 10125
rect -91 -2456 11101 6072
<< nwell >>
rect -200 10017 10450 10234
rect -200 -2250 115 10017
rect 10145 6344 10450 10017
rect 10246 6187 10450 6344
rect 5141 6186 10450 6187
rect 5141 5929 11210 6186
rect 9361 5860 11210 5929
rect 10895 -2250 11210 5860
rect -200 -2565 11210 -2250
<< mvpsubdiff >>
rect -322 10323 -262 10357
rect 10517 10323 10577 10357
rect -322 10297 -288 10323
rect 10543 10297 10577 10323
rect 10543 6313 10577 6344
rect 10543 6279 10615 6313
rect 11230 6279 11337 6313
rect 11303 6248 11337 6279
rect -322 -2656 -288 -2630
rect 11303 -2656 11337 -2630
rect -322 -2690 -262 -2656
rect 11277 -2690 11337 -2656
<< mvnsubdiff >>
rect -134 10148 10384 10168
rect -134 10114 -54 10148
rect 10304 10114 10384 10148
rect -134 10094 10384 10114
rect -134 10088 -60 10094
rect -134 -2419 -114 10088
rect -80 -2419 -60 10088
rect 10310 10088 10384 10094
rect 10310 6152 10330 10088
rect 10364 6152 10384 10088
rect 10310 6120 10384 6152
rect 10310 6101 11144 6120
rect 10310 6067 10364 6101
rect 11054 6072 11144 6101
rect 11054 6067 11090 6072
rect 10310 6046 11090 6067
rect -134 -2425 -60 -2419
rect 11070 -2410 11090 6046
rect 11124 -2410 11144 6072
rect 11070 -2425 11144 -2410
rect -134 -2445 11144 -2425
rect -134 -2479 -54 -2445
rect 11054 -2479 11144 -2445
rect -134 -2499 11144 -2479
<< mvpsubdiffcont >>
rect -262 10323 10517 10357
rect -322 -2630 -288 10297
rect 10543 6344 10577 10297
rect 10615 6279 11230 6313
rect 11303 -2630 11337 6248
rect -262 -2690 11277 -2656
<< mvnsubdiffcont >>
rect -54 10114 10304 10148
rect -114 -2419 -80 10088
rect 10330 6152 10364 10088
rect 10364 6067 11054 6101
rect 11090 -2410 11124 6072
rect -54 -2479 11054 -2445
<< locali >>
rect -322 10323 -262 10357
rect 10517 10323 10577 10357
rect -322 10317 10577 10323
rect -322 10297 -180 10317
rect -288 10268 -180 10297
rect 10415 10297 10577 10317
rect 10415 10268 10543 10297
rect -288 10235 10543 10268
rect -288 10154 -201 10235
rect -288 -2490 -276 10154
rect -224 -2490 -201 10154
rect 10449 10193 10543 10235
rect -114 10114 -54 10148
rect 10304 10114 10364 10148
rect -114 10088 10364 10114
rect -80 10065 10330 10088
rect -80 10015 84 10065
rect 10145 10015 10330 10065
rect -80 9970 10330 10015
rect -80 9936 63 9970
rect -80 -2285 -59 9936
rect -5 -2285 63 9936
rect 10175 9915 10330 9970
rect 10175 6151 10220 9915
rect 10272 6152 10330 9915
rect 10449 6344 10477 10193
rect 10534 6344 10543 10193
rect 12837 9463 12945 9473
rect 12837 9332 12850 9463
rect 12928 9332 12945 9463
rect 12837 9323 12945 9332
rect 12821 9011 12955 9026
rect 12821 8818 12834 9011
rect 12938 8818 12955 9011
rect 12821 8802 12955 8818
rect 11920 7236 12270 7248
rect 11920 7182 11945 7236
rect 12229 7182 12270 7236
rect 11920 7172 12270 7182
rect 10449 6313 10577 6344
rect 10449 6279 10615 6313
rect 11230 6279 11337 6313
rect 10449 6248 11337 6279
rect 10449 6186 11237 6248
rect 10272 6151 10364 6152
rect 10175 6067 10364 6151
rect 11054 6072 11124 6101
rect 11054 6067 11090 6072
rect 10175 6024 11090 6067
rect 10175 6008 10980 6024
rect 10175 5956 10226 6008
rect 10920 5956 10980 6008
rect 10175 5911 10980 5956
rect -80 -2290 63 -2285
rect 10934 -2290 10980 5911
rect -80 -2297 10980 -2290
rect 11036 -2297 11090 6024
rect -80 -2352 11090 -2297
rect -80 -2405 32 -2352
rect 10929 -2405 11090 -2352
rect -80 -2410 11090 -2405
rect -80 -2419 11124 -2410
rect -114 -2445 11124 -2419
rect -114 -2479 -54 -2445
rect 11054 -2479 11124 -2445
rect -288 -2566 -201 -2490
rect 11209 -2538 11237 6186
rect 11294 -2538 11303 6248
rect 11209 -2566 11303 -2538
rect -288 -2595 11303 -2566
rect -288 -2630 -153 -2595
rect -322 -2635 -153 -2630
rect 11184 -2630 11303 -2595
rect 11184 -2635 11337 -2630
rect -322 -2656 11337 -2635
rect -322 -2690 -262 -2656
rect 11277 -2690 11337 -2656
<< viali >>
rect -180 10268 10415 10317
rect -276 -2490 -224 10154
rect 84 10015 10145 10065
rect -59 -2285 -5 9936
rect 10220 6151 10272 9915
rect 10477 6344 10534 10193
rect 12850 9332 12928 9463
rect 12834 8818 12938 9011
rect 11945 7182 12229 7236
rect 10226 5956 10920 6008
rect 10980 -2297 11036 6024
rect 32 -2405 10929 -2352
rect 11237 -2538 11294 6248
rect -153 -2635 11184 -2595
<< metal1 >>
rect -322 10317 10577 10357
rect -322 10268 -180 10317
rect 10415 10268 10577 10317
rect -322 10235 10577 10268
rect -322 10154 -201 10235
rect -322 -2490 -276 10154
rect -224 -2490 -201 10154
rect 10449 10193 10577 10235
rect -72 10065 10290 10085
rect -72 10015 84 10065
rect 10145 10015 10290 10065
rect -72 10002 10290 10015
rect -72 9936 11 10002
rect 5161 9987 5347 10002
rect -72 -2285 -59 9936
rect -5 -2285 11 9936
rect 10207 9915 10290 10002
rect 3896 6109 3942 6237
rect 10207 6151 10220 9915
rect 10272 6151 10290 9915
rect 10449 7635 10477 10193
rect 10377 7627 10477 7635
rect 10534 9689 10577 10193
rect 10534 9688 11709 9689
rect 10534 9554 11726 9688
rect 10534 7627 10577 9554
rect 10549 6801 10577 7627
rect 11626 7192 11726 9554
rect 11920 7236 12270 7248
rect 11610 6801 11758 7192
rect 11920 7182 11945 7236
rect 12229 7182 12270 7236
rect 12363 7196 12523 9684
rect 12861 9473 12913 9873
rect 12837 9463 12945 9473
rect 12837 9332 12850 9463
rect 12928 9332 12945 9463
rect 12837 9323 12945 9332
rect 12861 9026 12913 9323
rect 12821 9011 12955 9026
rect 12821 8818 12834 9011
rect 12938 8818 12955 9011
rect 12821 8802 12955 8818
rect 11920 7174 12028 7182
rect 12200 7174 12270 7182
rect 11920 7172 12270 7174
rect 12028 7168 12200 7172
rect 12322 7130 12572 7196
rect 12322 6873 12336 7130
rect 12558 6873 12572 7130
rect 12322 6854 12572 6873
rect 12600 7147 12657 7213
rect 13166 7199 13266 9686
rect 12600 7137 12742 7147
rect 12600 6861 12639 7137
rect 12731 6861 12742 7137
rect 12600 6851 12742 6861
rect 13136 6801 13284 7199
rect 10549 6794 13284 6801
rect 10549 6564 11031 6794
rect 11327 6564 13284 6794
rect 10549 6558 13284 6564
rect 10549 6344 10577 6558
rect 12047 6417 12053 6420
rect 10377 6331 10577 6344
rect 10746 6371 12053 6417
rect 10207 6142 10290 6151
rect 10746 6109 10792 6371
rect 12047 6368 12053 6371
rect 12225 6368 12231 6420
rect 11137 6248 11337 6261
rect 97 6063 10792 6109
rect 10866 6164 11072 6175
rect 97 4054 143 6063
rect 10866 6027 10875 6164
rect 10207 6008 10875 6027
rect 10207 5956 10226 6008
rect 10207 5944 10875 5956
rect 11061 5944 11072 6164
rect 10866 5935 10980 5944
rect 97 4008 664 4054
rect -72 -2334 11 -2285
rect 10967 -2297 10980 5935
rect 11036 5935 11072 5944
rect 11036 -2297 11050 5935
rect 11309 5899 11337 6248
rect 11137 5891 11237 5899
rect 10967 -2334 11050 -2297
rect -72 -2352 11050 -2334
rect -72 -2405 32 -2352
rect 10929 -2405 11050 -2352
rect -72 -2417 11050 -2405
rect -322 -2520 -201 -2490
rect -322 -2566 3257 -2520
rect 11209 -2538 11237 5891
rect 11294 -2538 11337 5899
rect 11416 5843 11648 5852
rect 11416 5746 11422 5843
rect 11641 5746 11648 5843
rect 11416 3913 11648 5746
rect 11416 3425 11423 3913
rect 11639 3425 11648 3913
rect 11416 3413 11648 3425
rect 11209 -2566 11337 -2538
rect -322 -2595 11337 -2566
rect -322 -2635 -153 -2595
rect 11184 -2635 11337 -2595
rect -322 -2690 11337 -2635
rect -319 -2743 3257 -2690
<< via1 >>
rect 10377 6344 10477 7627
rect 10477 6344 10534 7627
rect 10534 6344 10549 7627
rect 12028 7182 12200 7226
rect 12028 7174 12200 7182
rect 12336 6873 12558 7130
rect 12639 6861 12731 7137
rect 11031 6564 11327 6794
rect 12053 6368 12225 6420
rect 10875 6024 11061 6164
rect 10875 6008 10980 6024
rect 10875 5956 10920 6008
rect 10920 5956 10980 6008
rect 10875 5944 10980 5956
rect 10980 5944 11036 6024
rect 11036 5944 11061 6024
rect 11137 5899 11237 6248
rect 11237 5899 11294 6248
rect 11294 5899 11309 6248
rect 11422 5746 11641 5843
rect 11423 3425 11639 3913
<< metal2 >>
rect 5161 9987 5347 10085
rect 10353 7627 10576 7653
rect 10353 6344 10377 7627
rect 10549 6450 10576 7627
rect 12022 7223 12028 7226
rect 12014 7177 12028 7223
rect 12022 7174 12028 7177
rect 12200 7174 12206 7226
rect 11026 6794 11336 6802
rect 11026 6564 11031 6794
rect 11327 6564 11336 6794
rect 11026 6450 11336 6564
rect 10549 6344 11336 6450
rect 12096 6426 12161 7174
rect 12318 7130 12569 7143
rect 12318 6873 12336 7130
rect 12558 6873 12569 7130
rect 12053 6420 12225 6426
rect 12053 6362 12225 6368
rect 4961 6175 5147 6257
rect 10355 6248 11336 6344
rect 10355 6227 11137 6248
rect 9712 6164 11072 6175
rect 9712 6163 10875 6164
rect 9712 5949 9725 6163
rect 10824 5949 10875 6163
rect 9712 5944 10875 5949
rect 11061 5944 11072 6164
rect 9712 5936 11072 5944
rect 9712 5935 11063 5936
rect 4961 5914 5147 5935
rect 11113 5899 11137 6227
rect 11309 5899 11336 6248
rect 12318 6164 12569 6873
rect 12318 5948 12331 6164
rect 12552 5948 12569 6164
rect 12318 5936 12569 5948
rect 12630 7137 12741 7146
rect 12630 6861 12639 7137
rect 12731 6861 12741 7137
rect 11113 4077 11336 5899
rect 12630 5849 12741 6861
rect 11413 5843 12741 5849
rect 11413 5746 11422 5843
rect 11641 5746 12741 5843
rect 11413 5738 12741 5746
rect 10640 3913 12121 3922
rect 10640 3425 11423 3913
rect 11639 3425 12121 3913
rect 10640 3417 12121 3425
rect -140 1871 198 1971
rect 10897 1738 11337 1838
rect -140 1636 198 1736
rect -140 1178 198 1278
<< via2 >>
rect 4961 5935 5147 6175
rect 9725 5949 10824 6163
rect 12331 5948 12552 6164
<< metal3 >>
rect 623 2142 723 7084
rect 1659 6114 1759 7545
rect 4954 6175 5158 6184
rect 835 6014 1759 6114
rect 2077 6160 4961 6175
rect 835 1343 935 6014
rect 2077 5948 2090 6160
rect 2488 5948 4961 6160
rect 2077 5935 4961 5948
rect 5147 6164 12571 6175
rect 5147 6163 12331 6164
rect 5147 5949 9725 6163
rect 10824 5949 12331 6163
rect 5147 5948 12331 5949
rect 12552 5948 12571 6164
rect 5147 5935 12571 5948
rect 4954 5927 5158 5935
<< via3 >>
rect 2090 5948 2488 6160
<< metal4 >>
rect 285 9775 1485 10036
rect 2570 9770 3770 10036
rect 285 6171 1485 6273
rect 2769 6216 6781 6936
rect 1685 6171 2501 6173
rect 285 6160 2501 6171
rect 285 5948 2090 6160
rect 2488 5948 2501 6160
rect 285 4660 2501 5948
rect 6061 5601 6781 6216
use cc_via2_3cut  cc_via2_3cut_0
timestamp 1717772055
transform 0 1 -639040 -1 0 518654
box 517199 639873 517310 640172
use cc_via2_3cut  cc_via2_3cut_1
timestamp 1717772055
transform 0 1 -639448 -1 0 519454
box 517199 639873 517310 640172
use comparator_bias  comparator_bias_0
timestamp 1721175533
transform -1 0 518254 0 1 -639855
box 508008 646042 518182 649916
use comparator_core_cload  comparator_core_cload_0
timestamp 1721179627
transform 1 0 -506133 0 1 -641069
box 506207 638825 517124 647001
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 0 1 11633 1 0 9302
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 0 -1 13261 -1 0 9494
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 0 -1 13261 -1 0 9686
box -66 -43 258 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 0 -1 13261 -1 0 9302
box -66 -43 2178 1671
<< labels >>
flabel metal2 -140 1871 198 1971 0 FreeSans 1600 0 0 0 VINP
port 1 nsew
flabel metal2 -140 1636 198 1736 0 FreeSans 1600 0 0 0 VINM
port 0 nsew
flabel metal4 285 9775 1485 10036 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal4 2570 9770 3770 10036 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal2 11113 4077 11336 5865 0 FreeSans 1600 270 0 0 DVSS
port 6 nsew
flabel metal2 10902 3417 11337 3922 0 FreeSans 1600 0 0 0 DVDD
port 5 nsew
flabel metal2 10911 1738 11337 1838 0 FreeSans 1200 0 0 0 VOUT
port 7 nsew
flabel metal2 -140 1178 198 1278 0 FreeSans 1600 0 0 0 CLOAD
port 8 nsew
flabel metal1 12861 9704 12913 9873 0 FreeSans 320 90 0 0 ENA
port 9 nsew
<< end >>
