magic
tech sky130A
magscale 1 2
timestamp 1717725805
<< error_p >>
rect -2069 598 2069 602
rect -2069 -530 -2039 598
rect -2003 532 2003 536
rect -2003 -464 -1973 532
rect 1973 -464 2003 532
rect 2039 -530 2069 598
<< nwell >>
rect -2039 -564 2039 598
<< mvpmos >>
rect -1945 -464 -1345 536
rect -1287 -464 -687 536
rect -629 -464 -29 536
rect 29 -464 629 536
rect 687 -464 1287 536
rect 1345 -464 1945 536
<< mvpdiff >>
rect -2003 524 -1945 536
rect -2003 -452 -1991 524
rect -1957 -452 -1945 524
rect -2003 -464 -1945 -452
rect -1345 524 -1287 536
rect -1345 -452 -1333 524
rect -1299 -452 -1287 524
rect -1345 -464 -1287 -452
rect -687 524 -629 536
rect -687 -452 -675 524
rect -641 -452 -629 524
rect -687 -464 -629 -452
rect -29 524 29 536
rect -29 -452 -17 524
rect 17 -452 29 524
rect -29 -464 29 -452
rect 629 524 687 536
rect 629 -452 641 524
rect 675 -452 687 524
rect 629 -464 687 -452
rect 1287 524 1345 536
rect 1287 -452 1299 524
rect 1333 -452 1345 524
rect 1287 -464 1345 -452
rect 1945 524 2003 536
rect 1945 -452 1957 524
rect 1991 -452 2003 524
rect 1945 -464 2003 -452
<< mvpdiffc >>
rect -1991 -452 -1957 524
rect -1333 -452 -1299 524
rect -675 -452 -641 524
rect -17 -452 17 524
rect 641 -452 675 524
rect 1299 -452 1333 524
rect 1957 -452 1991 524
<< poly >>
rect -1945 536 -1345 562
rect -1287 536 -687 562
rect -629 536 -29 562
rect 29 536 629 562
rect 687 536 1287 562
rect 1345 536 1945 562
rect -1945 -511 -1345 -464
rect -1945 -545 -1929 -511
rect -1361 -545 -1345 -511
rect -1945 -561 -1345 -545
rect -1287 -511 -687 -464
rect -1287 -545 -1271 -511
rect -703 -545 -687 -511
rect -1287 -561 -687 -545
rect -629 -511 -29 -464
rect -629 -545 -613 -511
rect -45 -545 -29 -511
rect -629 -561 -29 -545
rect 29 -511 629 -464
rect 29 -545 45 -511
rect 613 -545 629 -511
rect 29 -561 629 -545
rect 687 -511 1287 -464
rect 687 -545 703 -511
rect 1271 -545 1287 -511
rect 687 -561 1287 -545
rect 1345 -511 1945 -464
rect 1345 -545 1361 -511
rect 1929 -545 1945 -511
rect 1345 -561 1945 -545
<< polycont >>
rect -1929 -545 -1361 -511
rect -1271 -545 -703 -511
rect -613 -545 -45 -511
rect 45 -545 613 -511
rect 703 -545 1271 -511
rect 1361 -545 1929 -511
<< locali >>
rect -1991 524 -1957 540
rect -1991 -468 -1957 -452
rect -1333 524 -1299 540
rect -1333 -468 -1299 -452
rect -675 524 -641 540
rect -675 -468 -641 -452
rect -17 524 17 540
rect -17 -468 17 -452
rect 641 524 675 540
rect 641 -468 675 -452
rect 1299 524 1333 540
rect 1299 -468 1333 -452
rect 1957 524 1991 540
rect 1957 -468 1991 -452
rect -1945 -545 -1929 -511
rect -1361 -545 -1345 -511
rect -1287 -545 -1271 -511
rect -703 -545 -687 -511
rect -629 -545 -613 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 613 -545 629 -511
rect 687 -545 703 -511
rect 1271 -545 1287 -511
rect 1345 -545 1361 -511
rect 1929 -545 1945 -511
<< viali >>
rect -1991 -452 -1957 524
rect -1333 -452 -1299 524
rect -675 -452 -641 524
rect -17 -452 17 524
rect 641 -452 675 524
rect 1299 -452 1333 524
rect 1957 -452 1991 524
rect -1929 -545 -1361 -511
rect -1271 -545 -703 -511
rect -613 -545 -45 -511
rect 45 -545 613 -511
rect 703 -545 1271 -511
rect 1361 -545 1929 -511
<< metal1 >>
rect -1997 524 -1951 536
rect -1997 -452 -1991 524
rect -1957 -452 -1951 524
rect -1997 -464 -1951 -452
rect -1339 524 -1293 536
rect -1339 -452 -1333 524
rect -1299 -452 -1293 524
rect -1339 -464 -1293 -452
rect -681 524 -635 536
rect -681 -452 -675 524
rect -641 -452 -635 524
rect -681 -464 -635 -452
rect -23 524 23 536
rect -23 -452 -17 524
rect 17 -452 23 524
rect -23 -464 23 -452
rect 635 524 681 536
rect 635 -452 641 524
rect 675 -452 681 524
rect 635 -464 681 -452
rect 1293 524 1339 536
rect 1293 -452 1299 524
rect 1333 -452 1339 524
rect 1293 -464 1339 -452
rect 1951 524 1997 536
rect 1951 -452 1957 524
rect 1991 -452 1997 524
rect 1951 -464 1997 -452
rect -1941 -511 -1349 -505
rect -1941 -545 -1929 -511
rect -1361 -545 -1349 -511
rect -1941 -551 -1349 -545
rect -1283 -511 -691 -505
rect -1283 -545 -1271 -511
rect -703 -545 -691 -511
rect -1283 -551 -691 -545
rect -625 -511 -33 -505
rect -625 -545 -613 -511
rect -45 -545 -33 -511
rect -625 -551 -33 -545
rect 33 -511 625 -505
rect 33 -545 45 -511
rect 613 -545 625 -511
rect 33 -551 625 -545
rect 691 -511 1283 -505
rect 691 -545 703 -511
rect 1271 -545 1283 -511
rect 691 -551 1283 -545
rect 1349 -511 1941 -505
rect 1349 -545 1361 -511
rect 1929 -545 1941 -511
rect 1349 -551 1941 -545
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 3 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
