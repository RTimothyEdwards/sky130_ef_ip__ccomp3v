magic
tech sky130A
magscale 1 2
timestamp 1652806316
<< dnwell >>
rect -91 5652 10727 10125
rect -91 -156 9527 5652
<< nwell >>
rect -200 10017 10836 10234
rect -200 50 115 10017
rect 10521 6187 10836 10017
rect 5341 5929 10836 6187
rect 9361 5858 10836 5929
rect 9321 5543 10836 5858
rect 9321 50 9636 5543
rect -200 -265 9636 50
<< mvnsubdiff >>
rect -134 10148 10770 10168
rect -134 10114 -54 10148
rect 10690 10114 10770 10148
rect -134 10094 10770 10114
rect -134 10088 -60 10094
rect -134 -119 -114 10088
rect -80 -119 -60 10088
rect 10696 10088 10770 10094
rect 10696 5684 10716 10088
rect 10750 5684 10770 10088
rect 10696 5683 10770 5684
rect -134 -125 -60 -119
rect 9496 5663 10770 5683
rect 9496 5629 9594 5663
rect 10684 5629 10770 5663
rect 9496 5609 10770 5629
rect 9496 5575 9570 5609
rect 9496 -110 9516 5575
rect 9550 -110 9570 5575
rect 9496 -125 9570 -110
rect -134 -145 9570 -125
rect -134 -179 -54 -145
rect 9480 -179 9570 -145
rect -134 -199 9570 -179
<< mvnsubdiffcont >>
rect -54 10114 10690 10148
rect -114 -119 -80 10088
rect 10716 5684 10750 10088
rect 9594 5629 10684 5663
rect 9516 -110 9550 5575
rect -54 -179 9480 -145
<< locali >>
rect -114 10114 -54 10148
rect 10690 10114 10750 10148
rect -114 10088 10750 10114
rect -80 10065 10716 10088
rect -80 10015 84 10065
rect 10535 10015 10716 10065
rect -80 9970 10716 10015
rect -80 9936 63 9970
rect -80 15 -59 9936
rect -5 15 63 9936
rect 10565 9915 10716 9970
rect 10565 5851 10610 9915
rect 10662 5851 10716 9915
rect 10565 5833 10716 5851
rect -80 10 63 15
rect 9360 5785 10716 5833
rect 9360 5730 9501 5785
rect 10562 5730 10716 5785
rect 9360 5713 10716 5730
rect 9360 10 9406 5713
rect -80 3 9406 10
rect 9462 5684 10716 5713
rect 9462 5663 10750 5684
rect 9462 5629 9594 5663
rect 10684 5629 10750 5663
rect 9462 5575 9550 5629
rect 10565 5627 10730 5629
rect 9462 3 9516 5575
rect -80 -52 9516 3
rect -80 -105 32 -52
rect 9355 -105 9516 -52
rect -80 -110 9516 -105
rect 11025 3297 11082 3304
rect -80 -119 9550 -110
rect -114 -145 9550 -119
rect -114 -179 -54 -145
rect 9480 -179 9550 -145
<< viali >>
rect 84 10015 10535 10065
rect -59 15 -5 9936
rect 10610 5851 10662 9915
rect 9501 5730 10562 5785
rect 9406 3 9462 5713
rect 32 -105 9355 -52
rect 10233 3756 10532 3828
rect 11025 3174 11082 3297
<< metal1 >>
rect -72 10065 10680 10085
rect -72 10015 84 10065
rect 10535 10015 10680 10065
rect -72 10002 10680 10015
rect -72 9936 11 10002
rect 5161 9987 5347 10002
rect -72 15 -59 9936
rect -5 15 11 9936
rect 10597 9915 10680 10002
rect 10597 5851 10610 9915
rect 10662 5851 10680 9915
rect 10597 5798 10680 5851
rect -72 -34 11 15
rect 9393 5785 10680 5798
rect 9393 5730 9501 5785
rect 10562 5730 10680 5785
rect 9393 5715 10680 5730
rect 10739 6164 10990 6176
rect 10739 5944 10751 6164
rect 10977 5944 10990 6164
rect 9393 5713 9476 5715
rect 9393 3 9406 5713
rect 9462 3 9476 5713
rect 10739 5506 10990 5944
rect 10654 5410 10711 5421
rect 9911 438 10174 4739
rect 10654 4656 10711 4905
rect 10739 4673 10813 5506
rect 10841 4673 10887 5506
rect 10915 4673 10989 5506
rect 10378 4332 10444 4344
rect 10378 3840 10444 4148
rect 10208 3828 10549 3840
rect 10208 3756 10233 3828
rect 10532 3756 10549 3828
rect 10208 3745 10549 3756
rect 11019 3297 11088 3310
rect 11019 3174 11025 3297
rect 11082 3174 11088 3297
rect 11019 3096 11088 3174
rect 11019 2907 11088 2919
rect 11435 438 11698 4716
rect 9393 -34 9476 3
rect -72 -52 9476 -34
rect -72 -105 32 -52
rect 9355 -105 9476 -52
rect -72 -117 9476 -105
rect 9910 414 11698 438
rect 9910 121 9944 414
rect 11672 121 11698 414
rect 9910 -196 11698 121
<< via1 >>
rect 10751 5944 10977 6164
rect 10654 4905 10711 5410
rect 10378 4148 10444 4332
rect 11019 2919 11088 3096
rect 9944 121 11672 414
<< metal2 >>
rect 5161 9987 5347 10085
rect 5161 6175 5347 6257
rect 9712 6164 10990 6175
rect 9712 6163 10751 6164
rect 9712 5949 9725 6163
rect 10474 5949 10751 6163
rect 9712 5944 10751 5949
rect 10977 5944 10990 6164
rect 9712 5935 10990 5944
rect 5161 5914 5347 5935
rect 10636 4905 10654 5410
rect 10711 4905 11712 5410
rect 10371 4148 10378 4332
rect 10444 4227 10452 4332
rect 10444 4148 11765 4227
rect -24 3052 314 3152
rect 11012 3019 11019 3096
rect 9331 2919 11019 3019
rect 11088 2919 11097 3096
rect -24 2817 314 2917
rect 9910 414 11698 438
rect 9910 121 9944 414
rect 11672 121 11698 414
rect 9910 -196 11698 121
<< via2 >>
rect 5161 5935 5347 6175
rect 9725 5949 10474 6163
<< metal3 >>
rect 840 5782 900 6482
rect 1884 6137 1944 6464
rect 5154 6175 5358 6184
rect 1137 6077 1944 6137
rect 2077 6160 5161 6175
rect 1137 5787 1197 6077
rect 2077 5948 2090 6160
rect 2488 5948 5161 6160
rect 2077 5935 5161 5948
rect 5347 6163 10490 6175
rect 5347 5949 9725 6163
rect 10474 5949 10490 6163
rect 5347 5935 10490 5949
rect 5154 5927 5358 5935
<< via3 >>
rect 2090 5948 2488 6160
<< metal4 >>
rect 485 9775 1685 10036
rect 2770 9770 3970 10036
rect 485 6173 1685 6232
rect 485 6160 2501 6173
rect 485 5948 2090 6160
rect 2488 5948 2501 6160
rect 2769 6136 5221 6856
rect 485 5934 2501 5948
rect 485 5604 1685 5934
rect 4501 5601 5221 6136
use comparator_core  comparator_core_0
timestamp 1652806316
transform 1 0 -507679 0 1 -639888
box 507669 639956 517124 645817
use comparator_bias  comparator_bias_0
timestamp 1652806316
transform -1 0 518454 0 1 -639855
box 507806 646042 518382 649916
use sky130_fd_sc_hvl__lsbufhv2lv_1  sky130_fd_sc_hvl__lsbufhv2lv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1652806316
transform 0 1 10050 1 0 3048
box -66 -43 1698 1671
<< labels >>
flabel metal2 -24 2817 314 2917 0 FreeSans 1600 0 0 0 VINM
port 0 nsew
flabel metal2 -24 3052 314 3152 0 FreeSans 1600 0 0 0 VINP
port 1 nsew
flabel metal4 485 9775 1685 10036 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal4 2770 9770 3970 10036 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal2 11681 4148 11765 4227 0 FreeSans 1600 0 0 0 VOUT
port 4 nsew
flabel metal2 11277 4905 11712 5410 0 FreeSans 1600 0 0 0 DVDD
port 5 nsew
flabel metal2 9910 -196 11698 27 0 FreeSans 1600 0 0 0 DVSS
port 6 nsew
<< end >>
