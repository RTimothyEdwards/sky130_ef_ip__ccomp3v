magic
tech sky130A
magscale 1 2
timestamp 1717769301
<< checkpaint >>
rect 506138 644639 506205 644862
<< metal1 >>
rect 506138 644855 506205 644862
rect 506138 644639 506205 644646
<< via1 >>
rect 506138 644646 506205 644855
<< metal2 >>
rect 506138 644855 506205 644862
rect 506138 644639 506205 644646
<< end >>
