magic
tech sky130A
magscale 1 2
timestamp 1717725805
<< mvnmos >>
rect -1629 -531 -29 469
rect 29 -531 1629 469
<< mvndiff >>
rect -1687 457 -1629 469
rect -1687 -519 -1675 457
rect -1641 -519 -1629 457
rect -1687 -531 -1629 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 1629 457 1687 469
rect 1629 -519 1641 457
rect 1675 -519 1687 457
rect 1629 -531 1687 -519
<< mvndiffc >>
rect -1675 -519 -1641 457
rect -17 -519 17 457
rect 1641 -519 1675 457
<< poly >>
rect -1629 541 -29 557
rect -1629 507 -1613 541
rect -45 507 -29 541
rect -1629 469 -29 507
rect 29 541 1629 557
rect 29 507 45 541
rect 1613 507 1629 541
rect 29 469 1629 507
rect -1629 -557 -29 -531
rect 29 -557 1629 -531
<< polycont >>
rect -1613 507 -45 541
rect 45 507 1613 541
<< locali >>
rect -1629 507 -1613 541
rect -45 507 -29 541
rect 29 507 45 541
rect 1613 507 1629 541
rect -1675 457 -1641 473
rect -1675 -535 -1641 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 1641 457 1675 473
rect 1641 -535 1675 -519
<< viali >>
rect -1613 507 -45 541
rect 45 507 1613 541
rect -1675 -519 -1641 457
rect -17 -519 17 457
rect 1641 -519 1675 457
<< metal1 >>
rect -1625 541 -33 547
rect -1625 507 -1613 541
rect -45 507 -33 541
rect -1625 501 -33 507
rect 33 541 1625 547
rect 33 507 45 541
rect 1613 507 1625 541
rect 33 501 1625 507
rect -1681 457 -1635 469
rect -1681 -519 -1675 457
rect -1641 -519 -1635 457
rect -1681 -531 -1635 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 1635 457 1681 469
rect 1635 -519 1641 457
rect 1675 -519 1681 457
rect 1635 -531 1681 -519
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 8 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
