magic
tech sky130A
magscale 1 2
timestamp 1731000523
<< nwell >>
rect -358 -1415 358 1415
<< mvpmos >>
rect -100 118 100 1118
rect -100 -1118 100 -118
<< mvpdiff >>
rect -158 1106 -100 1118
rect -158 130 -146 1106
rect -112 130 -100 1106
rect -158 118 -100 130
rect 100 1106 158 1118
rect 100 130 112 1106
rect 146 130 158 1106
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -1106 -146 -130
rect -112 -1106 -100 -130
rect -158 -1118 -100 -1106
rect 100 -130 158 -118
rect 100 -1106 112 -130
rect 146 -1106 158 -130
rect 100 -1118 158 -1106
<< mvpdiffc >>
rect -146 130 -112 1106
rect 112 130 146 1106
rect -146 -1106 -112 -130
rect 112 -1106 146 -130
<< mvnsubdiff >>
rect -292 1337 292 1349
rect -292 1303 -184 1337
rect 184 1303 292 1337
rect -292 1291 292 1303
rect -292 1241 -234 1291
rect -292 -1241 -280 1241
rect -246 -1241 -234 1241
rect 234 1241 292 1291
rect -292 -1291 -234 -1241
rect 234 -1241 246 1241
rect 280 -1241 292 1241
rect 234 -1291 292 -1241
rect -292 -1303 292 -1291
rect -292 -1337 -184 -1303
rect 184 -1337 292 -1303
rect -292 -1349 292 -1337
<< mvnsubdiffcont >>
rect -184 1303 184 1337
rect -280 -1241 -246 1241
rect 246 -1241 280 1241
rect -184 -1337 184 -1303
<< poly >>
rect -100 1199 100 1215
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -100 1118 100 1165
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -1165 100 -1118
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -100 -1215 100 -1199
<< polycont >>
rect -84 1165 84 1199
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1199 84 -1165
<< locali >>
rect -280 1303 -184 1337
rect 184 1303 280 1337
rect -280 1241 -246 1303
rect 246 1241 280 1303
rect -100 1165 -84 1199
rect 84 1165 100 1199
rect -146 1106 -112 1122
rect -146 114 -112 130
rect 112 1106 146 1122
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -1122 -112 -1106
rect 112 -130 146 -114
rect 112 -1122 146 -1106
rect -100 -1199 -84 -1165
rect 84 -1199 100 -1165
rect -280 -1303 -246 -1241
rect 246 -1303 280 -1241
rect -280 -1337 -184 -1303
rect 184 -1337 280 -1303
<< viali >>
rect -84 1165 84 1199
rect -146 130 -112 1106
rect 112 130 146 1106
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1106 -112 -130
rect 112 -1106 146 -130
rect -84 -1199 84 -1165
<< metal1 >>
rect -96 1199 96 1205
rect -96 1165 -84 1199
rect 84 1165 96 1199
rect -96 1159 96 1165
rect -152 1106 -106 1118
rect -152 130 -146 1106
rect -112 130 -106 1106
rect -152 118 -106 130
rect 106 1106 152 1118
rect 106 130 112 1106
rect 146 130 152 1106
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -1106 -146 -130
rect -112 -1106 -106 -130
rect -152 -1118 -106 -1106
rect 106 -130 152 -118
rect 106 -1106 112 -130
rect 146 -1106 152 -130
rect 106 -1118 152 -1106
rect -96 -1165 96 -1159
rect -96 -1199 -84 -1165
rect 84 -1199 96 -1165
rect -96 -1205 96 -1199
<< properties >>
string FIXED_BBOX -263 -1320 263 1320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 1.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
