magic
tech sky130A
magscale 1 2
timestamp 1731019923
<< nwell >>
rect -458 -2297 458 2297
<< mvpmos >>
rect -200 -2000 200 2000
<< mvpdiff >>
rect -258 1988 -200 2000
rect -258 -1988 -246 1988
rect -212 -1988 -200 1988
rect -258 -2000 -200 -1988
rect 200 1988 258 2000
rect 200 -1988 212 1988
rect 246 -1988 258 1988
rect 200 -2000 258 -1988
<< mvpdiffc >>
rect -246 -1988 -212 1988
rect 212 -1988 246 1988
<< mvnsubdiff >>
rect -392 2219 392 2231
rect -392 2185 -284 2219
rect 284 2185 392 2219
rect -392 2173 392 2185
rect -392 2123 -334 2173
rect -392 -2123 -380 2123
rect -346 -2123 -334 2123
rect 334 2123 392 2173
rect -392 -2173 -334 -2123
rect 334 -2123 346 2123
rect 380 -2123 392 2123
rect 334 -2173 392 -2123
rect -392 -2185 392 -2173
rect -392 -2219 -284 -2185
rect 284 -2219 392 -2185
rect -392 -2231 392 -2219
<< mvnsubdiffcont >>
rect -284 2185 284 2219
rect -380 -2123 -346 2123
rect 346 -2123 380 2123
rect -284 -2219 284 -2185
<< poly >>
rect -200 2081 200 2097
rect -200 2047 -184 2081
rect 184 2047 200 2081
rect -200 2000 200 2047
rect -200 -2047 200 -2000
rect -200 -2081 -184 -2047
rect 184 -2081 200 -2047
rect -200 -2097 200 -2081
<< polycont >>
rect -184 2047 184 2081
rect -184 -2081 184 -2047
<< locali >>
rect -380 2185 -284 2219
rect 284 2185 380 2219
rect -380 2123 -346 2185
rect 346 2123 380 2185
rect -200 2047 -184 2081
rect 184 2047 200 2081
rect -246 1988 -212 2004
rect -246 -2004 -212 -1988
rect 212 1988 246 2004
rect 212 -2004 246 -1988
rect -200 -2081 -184 -2047
rect 184 -2081 200 -2047
rect -380 -2185 -346 -2123
rect 346 -2185 380 -2123
rect -380 -2219 -284 -2185
rect 284 -2219 380 -2185
<< viali >>
rect -184 2047 184 2081
rect -246 -1988 -212 1988
rect 212 -1988 246 1988
rect -184 -2081 184 -2047
<< metal1 >>
rect -196 2081 196 2087
rect -196 2047 -184 2081
rect 184 2047 196 2081
rect -196 2041 196 2047
rect -252 1988 -206 2000
rect -252 -1988 -246 1988
rect -212 -1988 -206 1988
rect -252 -2000 -206 -1988
rect 206 1988 252 2000
rect 206 -1988 212 1988
rect 246 -1988 252 1988
rect 206 -2000 252 -1988
rect -196 -2047 196 -2041
rect -196 -2081 -184 -2047
rect 184 -2081 196 -2047
rect -196 -2087 196 -2081
<< properties >>
string FIXED_BBOX -363 -2202 363 2202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 20.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
