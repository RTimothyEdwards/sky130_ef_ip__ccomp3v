magic
tech sky130A
magscale 1 2
timestamp 1731034391
<< dnwell >>
rect 52 304 8414 3984
rect 52 -3012 11076 304
<< nwell >>
rect -58 3778 8524 4094
rect -58 -2806 258 3778
rect 2532 3494 7612 3778
rect 2532 3392 4940 3494
rect 4172 3060 4940 3392
rect 4730 2314 4940 3060
rect 4778 324 4940 2314
rect 8208 414 8524 3778
rect 8208 98 11186 414
rect 10870 -2806 11186 98
rect -58 -3122 11186 -2806
<< mvnsubdiff >>
rect 9 4007 8443 4027
rect 9 3973 89 4007
rect 8328 3973 8443 4007
rect 9 3953 8443 3973
rect 9 3947 83 3953
rect 9 -2975 29 3947
rect 63 -2975 83 3947
rect 8369 3922 8443 3953
rect 8369 356 8389 3922
rect 8423 356 8443 3922
rect 8369 323 8443 356
rect 8369 303 11113 323
rect 8369 269 8482 303
rect 11000 269 11113 303
rect 8369 249 11113 269
rect 11039 220 11113 249
rect 9 -2981 83 -2975
rect 6346 -2981 6408 -2798
rect 11039 -2975 11059 220
rect 11093 -2975 11113 220
rect 11039 -2981 11113 -2975
rect 9 -3001 11113 -2981
rect 9 -3035 89 -3001
rect 11033 -3035 11113 -3001
rect 9 -3055 11113 -3035
<< mvnsubdiffcont >>
rect 89 3973 8328 4007
rect 29 -2975 63 3947
rect 8389 356 8423 3922
rect 8482 269 11000 303
rect 11059 -2975 11093 220
rect 89 -3035 11033 -3001
<< locali >>
rect 9 4013 8444 4028
rect 9 4007 108 4013
rect 8308 4007 8444 4013
rect 9 3973 89 4007
rect 8328 3973 8444 4007
rect 9 3967 108 3973
rect 8308 3967 8444 3973
rect 9 3953 8444 3967
rect 9 3947 84 3953
rect 9 3933 29 3947
rect 63 3933 84 3947
rect 9 -2947 23 3933
rect 65 -2947 84 3933
rect 8369 3922 8444 3953
rect 8369 3892 8389 3922
rect 8423 3892 8444 3922
rect 8369 387 8381 3892
rect 8426 387 8444 3892
rect 9215 3549 9413 3561
rect 9215 3434 9227 3549
rect 9399 3434 9413 3549
rect 9215 3423 9413 3434
rect 9218 2965 9399 2978
rect 9218 2844 9233 2965
rect 9386 2844 9399 2965
rect 9218 2833 9399 2844
rect 9890 1302 10224 1310
rect 9890 1202 10028 1302
rect 10206 1202 10224 1302
rect 9890 1192 10224 1202
rect 8369 356 8389 387
rect 8423 356 8444 387
rect 8369 324 8444 356
rect 8369 307 11114 324
rect 8369 305 10252 307
rect 8369 303 8497 305
rect 10068 303 10252 305
rect 10981 303 11114 307
rect 8369 269 8482 303
rect 11000 269 11114 303
rect 8369 262 8497 269
rect 10068 265 10252 269
rect 10981 265 11114 269
rect 10068 262 11114 265
rect 8369 249 11114 262
rect 11039 220 11114 249
rect 11039 195 11059 220
rect 11093 195 11114 220
rect 11039 -48 11052 195
rect 9 -2975 29 -2947
rect 63 -2975 84 -2947
rect 9 -2980 84 -2975
rect 6346 -2980 6408 -2798
rect 11038 -2951 11052 -48
rect 11096 -2951 11114 195
rect 11038 -2975 11059 -2951
rect 11093 -2975 11114 -2951
rect 11038 -2980 11114 -2975
rect 9 -2998 11114 -2980
rect 9 -3001 121 -2998
rect 11012 -3001 11114 -2998
rect 9 -3035 89 -3001
rect 11033 -3035 11114 -3001
rect 9 -3040 121 -3035
rect 11012 -3040 11114 -3035
rect 9 -3055 11114 -3040
<< viali >>
rect 108 4007 8308 4013
rect 108 3973 8308 4007
rect 108 3967 8308 3973
rect 23 -2947 29 3933
rect 29 -2947 63 3933
rect 63 -2947 65 3933
rect 8381 387 8389 3892
rect 8389 387 8423 3892
rect 8423 387 8426 3892
rect 9227 3434 9399 3549
rect 9233 2844 9386 2965
rect 10028 1202 10206 1302
rect 8497 303 10068 305
rect 10252 303 10981 307
rect 8497 269 10068 303
rect 10252 269 10981 303
rect 8497 262 10068 269
rect 10252 265 10981 269
rect 11052 -2951 11059 195
rect 11059 -2951 11093 195
rect 11093 -2951 11096 195
rect 121 -3001 11012 -2998
rect 121 -3035 11012 -3001
rect 121 -3040 11012 -3035
<< metal1 >>
rect 9 4013 8444 4028
rect 9 3967 108 4013
rect 8308 3967 8444 4013
rect 9 3953 8444 3967
rect 9 3933 84 3953
rect 9 3786 23 3933
rect -1 3776 23 3786
rect 65 3786 84 3933
rect 8369 3892 8444 3953
rect 65 3776 115 3786
rect 8369 3785 8381 3892
rect -1 3087 8 3776
rect 107 3087 115 3776
rect -1 3078 23 3087
rect 9 -2947 23 3078
rect 65 3078 115 3087
rect 8284 3770 8381 3785
rect 8426 3785 8444 3892
rect 9213 3808 9413 4008
rect 8426 3770 8473 3785
rect 8284 3089 8300 3770
rect 8456 3089 8473 3770
rect 8905 3402 9060 3586
rect 9286 3561 9338 3808
rect 9626 3692 9876 3704
rect 9215 3549 9413 3561
rect 9215 3434 9227 3549
rect 9399 3434 9413 3549
rect 9215 3423 9413 3434
rect 8284 3078 8381 3089
rect 65 -2947 84 3078
rect 8369 387 8381 3078
rect 8426 3078 8473 3089
rect 8426 387 8444 3078
rect 8906 1290 9060 3402
rect 9286 2978 9338 3423
rect 9626 3098 9634 3692
rect 9868 3098 9876 3692
rect 9626 3088 9876 3098
rect 9540 3012 9598 3028
rect 9218 2965 9399 2978
rect 9218 2844 9233 2965
rect 9386 2844 9399 2965
rect 9218 2833 9399 2844
rect 9286 2830 9338 2833
rect 9540 2792 9598 2806
rect 8906 1088 9062 1290
rect 9630 1284 9872 3088
rect 10010 1302 10344 1310
rect 10010 1202 10028 1302
rect 10206 1202 10344 1302
rect 10442 1292 10594 3586
rect 10010 1192 10344 1202
rect 8906 720 8912 1088
rect 9056 720 9062 1088
rect 8906 704 9062 720
rect 8369 324 8444 387
rect 8369 305 10096 324
rect 8369 262 8497 305
rect 10068 262 10096 305
rect 8369 249 10096 262
rect 10147 168 10182 1192
rect 10440 1098 10594 1292
rect 10322 1088 10594 1098
rect 10322 722 10328 1088
rect 10492 722 10594 1088
rect 10322 714 10594 722
rect 10232 307 11114 324
rect 10232 265 10252 307
rect 10981 265 11114 307
rect 10232 249 11114 265
rect 4792 134 10182 168
rect 11038 195 11114 249
rect 10736 -1268 10936 -1068
rect 10736 -1628 10936 -1428
rect 9 -2980 84 -2947
rect 6334 -2980 6420 -2821
rect 11038 -2951 11052 195
rect 11096 -2951 11114 195
rect 11038 -2980 11114 -2951
rect 9 -2998 11114 -2980
rect 9 -3040 121 -2998
rect 11012 -3040 11114 -2998
rect 9 -3055 11114 -3040
<< via1 >>
rect 8 3087 23 3776
rect 23 3087 65 3776
rect 65 3087 107 3776
rect 8300 3089 8381 3770
rect 8381 3089 8426 3770
rect 8426 3089 8456 3770
rect 9634 3098 9868 3692
rect 9540 2806 9598 3012
rect 8912 720 9056 1088
rect 10328 722 10492 1088
<< metal2 >>
rect -1 3776 10704 3786
rect -1 3087 8 3776
rect 107 3770 10704 3776
rect 107 3089 8300 3770
rect 8456 3692 10704 3770
rect 8456 3098 9634 3692
rect 9868 3098 10704 3692
rect 8456 3089 10704 3098
rect 107 3087 10704 3089
rect -1 3078 10704 3087
rect 8247 2806 9540 3012
rect 9598 2806 10704 3012
rect 10502 1736 10702 1792
rect 8046 1636 10702 1736
rect 10502 1592 10702 1636
rect 8288 1088 10704 1096
rect 8288 720 8912 1088
rect 9056 722 10328 1088
rect 10492 722 10704 1088
rect 9056 720 10704 722
rect 8288 714 10704 720
rect -13 -2786 6153 -2078
rect 6200 -2659 6555 -2077
rect 6199 -2787 6555 -2659
rect 6670 -2786 10764 -2658
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 0 1 8937 -1 0 3586
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1729530005
transform 0 -1 10565 1 0 3394
box -66 -43 258 897
use comparator_high_gain  x1
timestamp 1731033867
transform -1 0 11226 0 1 438
box 69 -3411 7124 3348
use scomp_bias  x2
timestamp 1731032193
transform -1 0 5269 0 1 -1439
box 323 -1349 5039 5225
use sky130_fd_sc_hvl__lsbuflv2hv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1731019923
transform 0 1 8937 -1 0 3394
box -66 -43 2178 1671
<< labels >>
flabel metal2 10502 1592 10702 1792 0 FreeSans 256 0 0 0 VOUT
port 0 nsew
flabel metal2 10500 2806 10700 3006 0 FreeSans 256 0 0 0 DVDD
port 1 nsew
flabel metal2 10482 3516 10682 3716 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal2 10504 808 10704 1008 0 FreeSans 256 0 0 0 DVSS
port 2 nsew
flabel metal1 10736 -1628 10936 -1428 0 FreeSans 256 0 0 0 VINM
port 6 nsew
flabel metal1 10736 -1268 10936 -1068 0 FreeSans 256 0 0 0 VINP
port 5 nsew
flabel metal2 6305 -2511 6505 -2311 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 9213 3808 9413 4008 0 FreeSans 256 0 0 0 ENA
port 7 nsew
<< end >>
